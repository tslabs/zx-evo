// bin2v output
// 

module bin2v(

	input  wire [15:0] in_addr,

	output reg  [ 7:0] out_word

);

	always @*
	case( in_addr )

		16'h0: out_word = 8'hF3;
		16'h1: out_word = 8'hAF;
		16'h2: out_word = 8'h11;
		16'h3: out_word = 8'hFF;
		16'h4: out_word = 8'hFF;
		16'h5: out_word = 8'hC3;
		16'h6: out_word = 8'hCB;
		16'h7: out_word = 8'h11;
		16'h8: out_word = 8'h2A;
		16'h9: out_word = 8'h5D;
		16'hA: out_word = 8'h5C;
		16'hB: out_word = 8'h22;
		16'hC: out_word = 8'h5F;
		16'hD: out_word = 8'h5C;
		16'hE: out_word = 8'h18;
		16'hF: out_word = 8'h43;
		16'h10: out_word = 8'hC3;
		16'h11: out_word = 8'hF2;
		16'h12: out_word = 8'h15;
		16'h13: out_word = 8'hFF;
		16'h14: out_word = 8'hFF;
		16'h15: out_word = 8'hFF;
		16'h16: out_word = 8'hFF;
		16'h17: out_word = 8'hFF;
		16'h18: out_word = 8'h2A;
		16'h19: out_word = 8'h5D;
		16'h1A: out_word = 8'h5C;
		16'h1B: out_word = 8'h7E;
		16'h1C: out_word = 8'hCD;
		16'h1D: out_word = 8'h7D;
		16'h1E: out_word = 8'h00;
		16'h1F: out_word = 8'hD0;
		16'h20: out_word = 8'hCD;
		16'h21: out_word = 8'h74;
		16'h22: out_word = 8'h00;
		16'h23: out_word = 8'h18;
		16'h24: out_word = 8'hF7;
		16'h25: out_word = 8'hFF;
		16'h26: out_word = 8'hFF;
		16'h27: out_word = 8'hFF;
		16'h28: out_word = 8'hC3;
		16'h29: out_word = 8'h5B;
		16'h2A: out_word = 8'h33;
		16'h2B: out_word = 8'hFF;
		16'h2C: out_word = 8'hFF;
		16'h2D: out_word = 8'hFF;
		16'h2E: out_word = 8'hFF;
		16'h2F: out_word = 8'hFF;
		16'h30: out_word = 8'hC5;
		16'h31: out_word = 8'h2A;
		16'h32: out_word = 8'h61;
		16'h33: out_word = 8'h5C;
		16'h34: out_word = 8'hE5;
		16'h35: out_word = 8'hC3;
		16'h36: out_word = 8'h9E;
		16'h37: out_word = 8'h16;
		16'h38: out_word = 8'hF5;
		16'h39: out_word = 8'hE5;
		16'h3A: out_word = 8'h2A;
		16'h3B: out_word = 8'h78;
		16'h3C: out_word = 8'h5C;
		16'h3D: out_word = 8'h23;
		16'h3E: out_word = 8'h22;
		16'h3F: out_word = 8'h78;
		16'h40: out_word = 8'h5C;
		16'h41: out_word = 8'h7C;
		16'h42: out_word = 8'hB5;
		16'h43: out_word = 8'h20;
		16'h44: out_word = 8'h03;
		16'h45: out_word = 8'hFD;
		16'h46: out_word = 8'h34;
		16'h47: out_word = 8'h40;
		16'h48: out_word = 8'hC5;
		16'h49: out_word = 8'hD5;
		16'h4A: out_word = 8'hCD;
		16'h4B: out_word = 8'h6E;
		16'h4C: out_word = 8'h38;
		16'h4D: out_word = 8'hD1;
		16'h4E: out_word = 8'hC1;
		16'h4F: out_word = 8'hE1;
		16'h50: out_word = 8'hF1;
		16'h51: out_word = 8'hFB;
		16'h52: out_word = 8'hC9;
		16'h53: out_word = 8'hE1;
		16'h54: out_word = 8'h6E;
		16'h55: out_word = 8'hFD;
		16'h56: out_word = 8'h75;
		16'h57: out_word = 8'h00;
		16'h58: out_word = 8'hED;
		16'h59: out_word = 8'h7B;
		16'h5A: out_word = 8'h3D;
		16'h5B: out_word = 8'h5C;
		16'h5C: out_word = 8'hC3;
		16'h5D: out_word = 8'hC5;
		16'h5E: out_word = 8'h16;
		16'h5F: out_word = 8'hFF;
		16'h60: out_word = 8'hFF;
		16'h61: out_word = 8'hFF;
		16'h62: out_word = 8'hFF;
		16'h63: out_word = 8'hFF;
		16'h64: out_word = 8'hFF;
		16'h65: out_word = 8'hFF;
		16'h66: out_word = 8'hF5;
		16'h67: out_word = 8'hE5;
		16'h68: out_word = 8'h2A;
		16'h69: out_word = 8'hB0;
		16'h6A: out_word = 8'h5C;
		16'h6B: out_word = 8'h7C;
		16'h6C: out_word = 8'hB5;
		16'h6D: out_word = 8'h20;
		16'h6E: out_word = 8'h01;
		16'h6F: out_word = 8'hE9;
		16'h70: out_word = 8'hE1;
		16'h71: out_word = 8'hF1;
		16'h72: out_word = 8'hED;
		16'h73: out_word = 8'h45;
		16'h74: out_word = 8'h2A;
		16'h75: out_word = 8'h5D;
		16'h76: out_word = 8'h5C;
		16'h77: out_word = 8'h23;
		16'h78: out_word = 8'h22;
		16'h79: out_word = 8'h5D;
		16'h7A: out_word = 8'h5C;
		16'h7B: out_word = 8'h7E;
		16'h7C: out_word = 8'hC9;
		16'h7D: out_word = 8'hFE;
		16'h7E: out_word = 8'h21;
		16'h7F: out_word = 8'hD0;
		16'h80: out_word = 8'hFE;
		16'h81: out_word = 8'h0D;
		16'h82: out_word = 8'hC8;
		16'h83: out_word = 8'hFE;
		16'h84: out_word = 8'h10;
		16'h85: out_word = 8'hD8;
		16'h86: out_word = 8'hFE;
		16'h87: out_word = 8'h18;
		16'h88: out_word = 8'h3F;
		16'h89: out_word = 8'hD8;
		16'h8A: out_word = 8'h23;
		16'h8B: out_word = 8'hFE;
		16'h8C: out_word = 8'h16;
		16'h8D: out_word = 8'h38;
		16'h8E: out_word = 8'h01;
		16'h8F: out_word = 8'h23;
		16'h90: out_word = 8'h37;
		16'h91: out_word = 8'h22;
		16'h92: out_word = 8'h5D;
		16'h93: out_word = 8'h5C;
		16'h94: out_word = 8'hC9;
		16'h95: out_word = 8'hBF;
		16'h96: out_word = 8'h52;
		16'h97: out_word = 8'h4E;
		16'h98: out_word = 8'hC4;
		16'h99: out_word = 8'h49;
		16'h9A: out_word = 8'h4E;
		16'h9B: out_word = 8'h4B;
		16'h9C: out_word = 8'h45;
		16'h9D: out_word = 8'h59;
		16'h9E: out_word = 8'hA4;
		16'h9F: out_word = 8'h50;
		16'hA0: out_word = 8'hC9;
		16'hA1: out_word = 8'h46;
		16'hA2: out_word = 8'hCE;
		16'hA3: out_word = 8'h50;
		16'hA4: out_word = 8'h4F;
		16'hA5: out_word = 8'h49;
		16'hA6: out_word = 8'h4E;
		16'hA7: out_word = 8'hD4;
		16'hA8: out_word = 8'h53;
		16'hA9: out_word = 8'h43;
		16'hAA: out_word = 8'h52;
		16'hAB: out_word = 8'h45;
		16'hAC: out_word = 8'h45;
		16'hAD: out_word = 8'h4E;
		16'hAE: out_word = 8'hA4;
		16'hAF: out_word = 8'h41;
		16'hB0: out_word = 8'h54;
		16'hB1: out_word = 8'h54;
		16'hB2: out_word = 8'hD2;
		16'hB3: out_word = 8'h41;
		16'hB4: out_word = 8'hD4;
		16'hB5: out_word = 8'h54;
		16'hB6: out_word = 8'h41;
		16'hB7: out_word = 8'hC2;
		16'hB8: out_word = 8'h56;
		16'hB9: out_word = 8'h41;
		16'hBA: out_word = 8'h4C;
		16'hBB: out_word = 8'hA4;
		16'hBC: out_word = 8'h43;
		16'hBD: out_word = 8'h4F;
		16'hBE: out_word = 8'h44;
		16'hBF: out_word = 8'hC5;
		16'hC0: out_word = 8'h56;
		16'hC1: out_word = 8'h41;
		16'hC2: out_word = 8'hCC;
		16'hC3: out_word = 8'h4C;
		16'hC4: out_word = 8'h45;
		16'hC5: out_word = 8'hCE;
		16'hC6: out_word = 8'h53;
		16'hC7: out_word = 8'h49;
		16'hC8: out_word = 8'hCE;
		16'hC9: out_word = 8'h43;
		16'hCA: out_word = 8'h4F;
		16'hCB: out_word = 8'hD3;
		16'hCC: out_word = 8'h54;
		16'hCD: out_word = 8'h41;
		16'hCE: out_word = 8'hCE;
		16'hCF: out_word = 8'h41;
		16'hD0: out_word = 8'h53;
		16'hD1: out_word = 8'hCE;
		16'hD2: out_word = 8'h41;
		16'hD3: out_word = 8'h43;
		16'hD4: out_word = 8'hD3;
		16'hD5: out_word = 8'h41;
		16'hD6: out_word = 8'h54;
		16'hD7: out_word = 8'hCE;
		16'hD8: out_word = 8'h4C;
		16'hD9: out_word = 8'hCE;
		16'hDA: out_word = 8'h45;
		16'hDB: out_word = 8'h58;
		16'hDC: out_word = 8'hD0;
		16'hDD: out_word = 8'h49;
		16'hDE: out_word = 8'h4E;
		16'hDF: out_word = 8'hD4;
		16'hE0: out_word = 8'h53;
		16'hE1: out_word = 8'h51;
		16'hE2: out_word = 8'hD2;
		16'hE3: out_word = 8'h53;
		16'hE4: out_word = 8'h47;
		16'hE5: out_word = 8'hCE;
		16'hE6: out_word = 8'h41;
		16'hE7: out_word = 8'h42;
		16'hE8: out_word = 8'hD3;
		16'hE9: out_word = 8'h50;
		16'hEA: out_word = 8'h45;
		16'hEB: out_word = 8'h45;
		16'hEC: out_word = 8'hCB;
		16'hED: out_word = 8'h49;
		16'hEE: out_word = 8'hCE;
		16'hEF: out_word = 8'h55;
		16'hF0: out_word = 8'h53;
		16'hF1: out_word = 8'hD2;
		16'hF2: out_word = 8'h53;
		16'hF3: out_word = 8'h54;
		16'hF4: out_word = 8'h52;
		16'hF5: out_word = 8'hA4;
		16'hF6: out_word = 8'h43;
		16'hF7: out_word = 8'h48;
		16'hF8: out_word = 8'h52;
		16'hF9: out_word = 8'hA4;
		16'hFA: out_word = 8'h4E;
		16'hFB: out_word = 8'h4F;
		16'hFC: out_word = 8'hD4;
		16'hFD: out_word = 8'h42;
		16'hFE: out_word = 8'h49;
		16'hFF: out_word = 8'hCE;
		16'h100: out_word = 8'h4F;
		16'h101: out_word = 8'hD2;
		16'h102: out_word = 8'h41;
		16'h103: out_word = 8'h4E;
		16'h104: out_word = 8'hC4;
		16'h105: out_word = 8'h3C;
		16'h106: out_word = 8'hBD;
		16'h107: out_word = 8'h3E;
		16'h108: out_word = 8'hBD;
		16'h109: out_word = 8'h3C;
		16'h10A: out_word = 8'hBE;
		16'h10B: out_word = 8'h4C;
		16'h10C: out_word = 8'h49;
		16'h10D: out_word = 8'h4E;
		16'h10E: out_word = 8'hC5;
		16'h10F: out_word = 8'h54;
		16'h110: out_word = 8'h48;
		16'h111: out_word = 8'h45;
		16'h112: out_word = 8'hCE;
		16'h113: out_word = 8'h54;
		16'h114: out_word = 8'hCF;
		16'h115: out_word = 8'h53;
		16'h116: out_word = 8'h54;
		16'h117: out_word = 8'h45;
		16'h118: out_word = 8'hD0;
		16'h119: out_word = 8'h44;
		16'h11A: out_word = 8'h45;
		16'h11B: out_word = 8'h46;
		16'h11C: out_word = 8'h20;
		16'h11D: out_word = 8'h46;
		16'h11E: out_word = 8'hCE;
		16'h11F: out_word = 8'h43;
		16'h120: out_word = 8'h41;
		16'h121: out_word = 8'hD4;
		16'h122: out_word = 8'h46;
		16'h123: out_word = 8'h4F;
		16'h124: out_word = 8'h52;
		16'h125: out_word = 8'h4D;
		16'h126: out_word = 8'h41;
		16'h127: out_word = 8'hD4;
		16'h128: out_word = 8'h4D;
		16'h129: out_word = 8'h4F;
		16'h12A: out_word = 8'h56;
		16'h12B: out_word = 8'hC5;
		16'h12C: out_word = 8'h45;
		16'h12D: out_word = 8'h52;
		16'h12E: out_word = 8'h41;
		16'h12F: out_word = 8'h53;
		16'h130: out_word = 8'hC5;
		16'h131: out_word = 8'h4F;
		16'h132: out_word = 8'h50;
		16'h133: out_word = 8'h45;
		16'h134: out_word = 8'h4E;
		16'h135: out_word = 8'h20;
		16'h136: out_word = 8'hA3;
		16'h137: out_word = 8'h43;
		16'h138: out_word = 8'h4C;
		16'h139: out_word = 8'h4F;
		16'h13A: out_word = 8'h53;
		16'h13B: out_word = 8'h45;
		16'h13C: out_word = 8'h20;
		16'h13D: out_word = 8'hA3;
		16'h13E: out_word = 8'h4D;
		16'h13F: out_word = 8'h45;
		16'h140: out_word = 8'h52;
		16'h141: out_word = 8'h47;
		16'h142: out_word = 8'hC5;
		16'h143: out_word = 8'h56;
		16'h144: out_word = 8'h45;
		16'h145: out_word = 8'h52;
		16'h146: out_word = 8'h49;
		16'h147: out_word = 8'h46;
		16'h148: out_word = 8'hD9;
		16'h149: out_word = 8'h42;
		16'h14A: out_word = 8'h45;
		16'h14B: out_word = 8'h45;
		16'h14C: out_word = 8'hD0;
		16'h14D: out_word = 8'h43;
		16'h14E: out_word = 8'h49;
		16'h14F: out_word = 8'h52;
		16'h150: out_word = 8'h43;
		16'h151: out_word = 8'h4C;
		16'h152: out_word = 8'hC5;
		16'h153: out_word = 8'h49;
		16'h154: out_word = 8'h4E;
		16'h155: out_word = 8'hCB;
		16'h156: out_word = 8'h50;
		16'h157: out_word = 8'h41;
		16'h158: out_word = 8'h50;
		16'h159: out_word = 8'h45;
		16'h15A: out_word = 8'hD2;
		16'h15B: out_word = 8'h46;
		16'h15C: out_word = 8'h4C;
		16'h15D: out_word = 8'h41;
		16'h15E: out_word = 8'h53;
		16'h15F: out_word = 8'hC8;
		16'h160: out_word = 8'h42;
		16'h161: out_word = 8'h52;
		16'h162: out_word = 8'h49;
		16'h163: out_word = 8'h47;
		16'h164: out_word = 8'h48;
		16'h165: out_word = 8'hD4;
		16'h166: out_word = 8'h49;
		16'h167: out_word = 8'h4E;
		16'h168: out_word = 8'h56;
		16'h169: out_word = 8'h45;
		16'h16A: out_word = 8'h52;
		16'h16B: out_word = 8'h53;
		16'h16C: out_word = 8'hC5;
		16'h16D: out_word = 8'h4F;
		16'h16E: out_word = 8'h56;
		16'h16F: out_word = 8'h45;
		16'h170: out_word = 8'hD2;
		16'h171: out_word = 8'h4F;
		16'h172: out_word = 8'h55;
		16'h173: out_word = 8'hD4;
		16'h174: out_word = 8'h4C;
		16'h175: out_word = 8'h50;
		16'h176: out_word = 8'h52;
		16'h177: out_word = 8'h49;
		16'h178: out_word = 8'h4E;
		16'h179: out_word = 8'hD4;
		16'h17A: out_word = 8'h4C;
		16'h17B: out_word = 8'h4C;
		16'h17C: out_word = 8'h49;
		16'h17D: out_word = 8'h53;
		16'h17E: out_word = 8'hD4;
		16'h17F: out_word = 8'h53;
		16'h180: out_word = 8'h54;
		16'h181: out_word = 8'h4F;
		16'h182: out_word = 8'hD0;
		16'h183: out_word = 8'h52;
		16'h184: out_word = 8'h45;
		16'h185: out_word = 8'h41;
		16'h186: out_word = 8'hC4;
		16'h187: out_word = 8'h44;
		16'h188: out_word = 8'h41;
		16'h189: out_word = 8'h54;
		16'h18A: out_word = 8'hC1;
		16'h18B: out_word = 8'h52;
		16'h18C: out_word = 8'h45;
		16'h18D: out_word = 8'h53;
		16'h18E: out_word = 8'h54;
		16'h18F: out_word = 8'h4F;
		16'h190: out_word = 8'h52;
		16'h191: out_word = 8'hC5;
		16'h192: out_word = 8'h4E;
		16'h193: out_word = 8'h45;
		16'h194: out_word = 8'hD7;
		16'h195: out_word = 8'h42;
		16'h196: out_word = 8'h4F;
		16'h197: out_word = 8'h52;
		16'h198: out_word = 8'h44;
		16'h199: out_word = 8'h45;
		16'h19A: out_word = 8'hD2;
		16'h19B: out_word = 8'h43;
		16'h19C: out_word = 8'h4F;
		16'h19D: out_word = 8'h4E;
		16'h19E: out_word = 8'h54;
		16'h19F: out_word = 8'h49;
		16'h1A0: out_word = 8'h4E;
		16'h1A1: out_word = 8'h55;
		16'h1A2: out_word = 8'hC5;
		16'h1A3: out_word = 8'h44;
		16'h1A4: out_word = 8'h49;
		16'h1A5: out_word = 8'hCD;
		16'h1A6: out_word = 8'h52;
		16'h1A7: out_word = 8'h45;
		16'h1A8: out_word = 8'hCD;
		16'h1A9: out_word = 8'h46;
		16'h1AA: out_word = 8'h4F;
		16'h1AB: out_word = 8'hD2;
		16'h1AC: out_word = 8'h47;
		16'h1AD: out_word = 8'h4F;
		16'h1AE: out_word = 8'h20;
		16'h1AF: out_word = 8'h54;
		16'h1B0: out_word = 8'hCF;
		16'h1B1: out_word = 8'h47;
		16'h1B2: out_word = 8'h4F;
		16'h1B3: out_word = 8'h20;
		16'h1B4: out_word = 8'h53;
		16'h1B5: out_word = 8'h55;
		16'h1B6: out_word = 8'hC2;
		16'h1B7: out_word = 8'h49;
		16'h1B8: out_word = 8'h4E;
		16'h1B9: out_word = 8'h50;
		16'h1BA: out_word = 8'h55;
		16'h1BB: out_word = 8'hD4;
		16'h1BC: out_word = 8'h4C;
		16'h1BD: out_word = 8'h4F;
		16'h1BE: out_word = 8'h41;
		16'h1BF: out_word = 8'hC4;
		16'h1C0: out_word = 8'h4C;
		16'h1C1: out_word = 8'h49;
		16'h1C2: out_word = 8'h53;
		16'h1C3: out_word = 8'hD4;
		16'h1C4: out_word = 8'h4C;
		16'h1C5: out_word = 8'h45;
		16'h1C6: out_word = 8'hD4;
		16'h1C7: out_word = 8'h50;
		16'h1C8: out_word = 8'h41;
		16'h1C9: out_word = 8'h55;
		16'h1CA: out_word = 8'h53;
		16'h1CB: out_word = 8'hC5;
		16'h1CC: out_word = 8'h4E;
		16'h1CD: out_word = 8'h45;
		16'h1CE: out_word = 8'h58;
		16'h1CF: out_word = 8'hD4;
		16'h1D0: out_word = 8'h50;
		16'h1D1: out_word = 8'h4F;
		16'h1D2: out_word = 8'h4B;
		16'h1D3: out_word = 8'hC5;
		16'h1D4: out_word = 8'h50;
		16'h1D5: out_word = 8'h52;
		16'h1D6: out_word = 8'h49;
		16'h1D7: out_word = 8'h4E;
		16'h1D8: out_word = 8'hD4;
		16'h1D9: out_word = 8'h50;
		16'h1DA: out_word = 8'h4C;
		16'h1DB: out_word = 8'h4F;
		16'h1DC: out_word = 8'hD4;
		16'h1DD: out_word = 8'h52;
		16'h1DE: out_word = 8'h55;
		16'h1DF: out_word = 8'hCE;
		16'h1E0: out_word = 8'h53;
		16'h1E1: out_word = 8'h41;
		16'h1E2: out_word = 8'h56;
		16'h1E3: out_word = 8'hC5;
		16'h1E4: out_word = 8'h52;
		16'h1E5: out_word = 8'h41;
		16'h1E6: out_word = 8'h4E;
		16'h1E7: out_word = 8'h44;
		16'h1E8: out_word = 8'h4F;
		16'h1E9: out_word = 8'h4D;
		16'h1EA: out_word = 8'h49;
		16'h1EB: out_word = 8'h5A;
		16'h1EC: out_word = 8'hC5;
		16'h1ED: out_word = 8'h49;
		16'h1EE: out_word = 8'hC6;
		16'h1EF: out_word = 8'h43;
		16'h1F0: out_word = 8'h4C;
		16'h1F1: out_word = 8'hD3;
		16'h1F2: out_word = 8'h44;
		16'h1F3: out_word = 8'h52;
		16'h1F4: out_word = 8'h41;
		16'h1F5: out_word = 8'hD7;
		16'h1F6: out_word = 8'h43;
		16'h1F7: out_word = 8'h4C;
		16'h1F8: out_word = 8'h45;
		16'h1F9: out_word = 8'h41;
		16'h1FA: out_word = 8'hD2;
		16'h1FB: out_word = 8'h52;
		16'h1FC: out_word = 8'h45;
		16'h1FD: out_word = 8'h54;
		16'h1FE: out_word = 8'h55;
		16'h1FF: out_word = 8'h52;
		16'h200: out_word = 8'hCE;
		16'h201: out_word = 8'h43;
		16'h202: out_word = 8'h4F;
		16'h203: out_word = 8'h50;
		16'h204: out_word = 8'hD9;
		16'h205: out_word = 8'h42;
		16'h206: out_word = 8'h48;
		16'h207: out_word = 8'h59;
		16'h208: out_word = 8'h36;
		16'h209: out_word = 8'h35;
		16'h20A: out_word = 8'h54;
		16'h20B: out_word = 8'h47;
		16'h20C: out_word = 8'h56;
		16'h20D: out_word = 8'h4E;
		16'h20E: out_word = 8'h4A;
		16'h20F: out_word = 8'h55;
		16'h210: out_word = 8'h37;
		16'h211: out_word = 8'h34;
		16'h212: out_word = 8'h52;
		16'h213: out_word = 8'h46;
		16'h214: out_word = 8'h43;
		16'h215: out_word = 8'h4D;
		16'h216: out_word = 8'h4B;
		16'h217: out_word = 8'h49;
		16'h218: out_word = 8'h38;
		16'h219: out_word = 8'h33;
		16'h21A: out_word = 8'h45;
		16'h21B: out_word = 8'h44;
		16'h21C: out_word = 8'h58;
		16'h21D: out_word = 8'h0E;
		16'h21E: out_word = 8'h4C;
		16'h21F: out_word = 8'h4F;
		16'h220: out_word = 8'h39;
		16'h221: out_word = 8'h32;
		16'h222: out_word = 8'h57;
		16'h223: out_word = 8'h53;
		16'h224: out_word = 8'h5A;
		16'h225: out_word = 8'h20;
		16'h226: out_word = 8'h0D;
		16'h227: out_word = 8'h50;
		16'h228: out_word = 8'h30;
		16'h229: out_word = 8'h31;
		16'h22A: out_word = 8'h51;
		16'h22B: out_word = 8'h41;
		16'h22C: out_word = 8'hE3;
		16'h22D: out_word = 8'hC4;
		16'h22E: out_word = 8'hE0;
		16'h22F: out_word = 8'hE4;
		16'h230: out_word = 8'hB4;
		16'h231: out_word = 8'hBC;
		16'h232: out_word = 8'hBD;
		16'h233: out_word = 8'hBB;
		16'h234: out_word = 8'hAF;
		16'h235: out_word = 8'hB0;
		16'h236: out_word = 8'hB1;
		16'h237: out_word = 8'hC0;
		16'h238: out_word = 8'hA7;
		16'h239: out_word = 8'hA6;
		16'h23A: out_word = 8'hBE;
		16'h23B: out_word = 8'hAD;
		16'h23C: out_word = 8'hB2;
		16'h23D: out_word = 8'hBA;
		16'h23E: out_word = 8'hE5;
		16'h23F: out_word = 8'hA5;
		16'h240: out_word = 8'hC2;
		16'h241: out_word = 8'hE1;
		16'h242: out_word = 8'hB3;
		16'h243: out_word = 8'hB9;
		16'h244: out_word = 8'hC1;
		16'h245: out_word = 8'hB8;
		16'h246: out_word = 8'h7E;
		16'h247: out_word = 8'hDC;
		16'h248: out_word = 8'hDA;
		16'h249: out_word = 8'h5C;
		16'h24A: out_word = 8'hB7;
		16'h24B: out_word = 8'h7B;
		16'h24C: out_word = 8'h7D;
		16'h24D: out_word = 8'hD8;
		16'h24E: out_word = 8'hBF;
		16'h24F: out_word = 8'hAE;
		16'h250: out_word = 8'hAA;
		16'h251: out_word = 8'hAB;
		16'h252: out_word = 8'hDD;
		16'h253: out_word = 8'hDE;
		16'h254: out_word = 8'hDF;
		16'h255: out_word = 8'h7F;
		16'h256: out_word = 8'hB5;
		16'h257: out_word = 8'hD6;
		16'h258: out_word = 8'h7C;
		16'h259: out_word = 8'hD5;
		16'h25A: out_word = 8'h5D;
		16'h25B: out_word = 8'hDB;
		16'h25C: out_word = 8'hB6;
		16'h25D: out_word = 8'hD9;
		16'h25E: out_word = 8'h5B;
		16'h25F: out_word = 8'hD7;
		16'h260: out_word = 8'h0C;
		16'h261: out_word = 8'h07;
		16'h262: out_word = 8'h06;
		16'h263: out_word = 8'h04;
		16'h264: out_word = 8'h05;
		16'h265: out_word = 8'h08;
		16'h266: out_word = 8'h0A;
		16'h267: out_word = 8'h0B;
		16'h268: out_word = 8'h09;
		16'h269: out_word = 8'h0F;
		16'h26A: out_word = 8'hE2;
		16'h26B: out_word = 8'h2A;
		16'h26C: out_word = 8'h3F;
		16'h26D: out_word = 8'hCD;
		16'h26E: out_word = 8'hC8;
		16'h26F: out_word = 8'hCC;
		16'h270: out_word = 8'hCB;
		16'h271: out_word = 8'h5E;
		16'h272: out_word = 8'hAC;
		16'h273: out_word = 8'h2D;
		16'h274: out_word = 8'h2B;
		16'h275: out_word = 8'h3D;
		16'h276: out_word = 8'h2E;
		16'h277: out_word = 8'h2C;
		16'h278: out_word = 8'h3B;
		16'h279: out_word = 8'h22;
		16'h27A: out_word = 8'hC7;
		16'h27B: out_word = 8'h3C;
		16'h27C: out_word = 8'hC3;
		16'h27D: out_word = 8'h3E;
		16'h27E: out_word = 8'hC5;
		16'h27F: out_word = 8'h2F;
		16'h280: out_word = 8'hC9;
		16'h281: out_word = 8'h60;
		16'h282: out_word = 8'hC6;
		16'h283: out_word = 8'h3A;
		16'h284: out_word = 8'hD0;
		16'h285: out_word = 8'hCE;
		16'h286: out_word = 8'hA8;
		16'h287: out_word = 8'hCA;
		16'h288: out_word = 8'hD3;
		16'h289: out_word = 8'hD4;
		16'h28A: out_word = 8'hD1;
		16'h28B: out_word = 8'hD2;
		16'h28C: out_word = 8'hA9;
		16'h28D: out_word = 8'hCF;
		16'h28E: out_word = 8'h2E;
		16'h28F: out_word = 8'h2F;
		16'h290: out_word = 8'h11;
		16'h291: out_word = 8'hFF;
		16'h292: out_word = 8'hFF;
		16'h293: out_word = 8'h01;
		16'h294: out_word = 8'hFE;
		16'h295: out_word = 8'hFE;
		16'h296: out_word = 8'hED;
		16'h297: out_word = 8'h78;
		16'h298: out_word = 8'h2F;
		16'h299: out_word = 8'hE6;
		16'h29A: out_word = 8'h1F;
		16'h29B: out_word = 8'h28;
		16'h29C: out_word = 8'h0E;
		16'h29D: out_word = 8'h67;
		16'h29E: out_word = 8'h7D;
		16'h29F: out_word = 8'h14;
		16'h2A0: out_word = 8'hC0;
		16'h2A1: out_word = 8'hD6;
		16'h2A2: out_word = 8'h08;
		16'h2A3: out_word = 8'hCB;
		16'h2A4: out_word = 8'h3C;
		16'h2A5: out_word = 8'h30;
		16'h2A6: out_word = 8'hFA;
		16'h2A7: out_word = 8'h53;
		16'h2A8: out_word = 8'h5F;
		16'h2A9: out_word = 8'h20;
		16'h2AA: out_word = 8'hF4;
		16'h2AB: out_word = 8'h2D;
		16'h2AC: out_word = 8'hCB;
		16'h2AD: out_word = 8'h00;
		16'h2AE: out_word = 8'h38;
		16'h2AF: out_word = 8'hE6;
		16'h2B0: out_word = 8'h7A;
		16'h2B1: out_word = 8'h3C;
		16'h2B2: out_word = 8'hC8;
		16'h2B3: out_word = 8'hFE;
		16'h2B4: out_word = 8'h28;
		16'h2B5: out_word = 8'hC8;
		16'h2B6: out_word = 8'hFE;
		16'h2B7: out_word = 8'h19;
		16'h2B8: out_word = 8'hC8;
		16'h2B9: out_word = 8'h7B;
		16'h2BA: out_word = 8'h5A;
		16'h2BB: out_word = 8'h57;
		16'h2BC: out_word = 8'hFE;
		16'h2BD: out_word = 8'h18;
		16'h2BE: out_word = 8'hC9;
		16'h2BF: out_word = 8'hCD;
		16'h2C0: out_word = 8'h8E;
		16'h2C1: out_word = 8'h02;
		16'h2C2: out_word = 8'hC0;
		16'h2C3: out_word = 8'h21;
		16'h2C4: out_word = 8'h00;
		16'h2C5: out_word = 8'h5C;
		16'h2C6: out_word = 8'hCB;
		16'h2C7: out_word = 8'h7E;
		16'h2C8: out_word = 8'h20;
		16'h2C9: out_word = 8'h07;
		16'h2CA: out_word = 8'h23;
		16'h2CB: out_word = 8'h35;
		16'h2CC: out_word = 8'h2B;
		16'h2CD: out_word = 8'h20;
		16'h2CE: out_word = 8'h02;
		16'h2CF: out_word = 8'h36;
		16'h2D0: out_word = 8'hFF;
		16'h2D1: out_word = 8'h7D;
		16'h2D2: out_word = 8'h21;
		16'h2D3: out_word = 8'h04;
		16'h2D4: out_word = 8'h5C;
		16'h2D5: out_word = 8'hBD;
		16'h2D6: out_word = 8'h20;
		16'h2D7: out_word = 8'hEE;
		16'h2D8: out_word = 8'hCD;
		16'h2D9: out_word = 8'h1E;
		16'h2DA: out_word = 8'h03;
		16'h2DB: out_word = 8'hD0;
		16'h2DC: out_word = 8'h21;
		16'h2DD: out_word = 8'h00;
		16'h2DE: out_word = 8'h5C;
		16'h2DF: out_word = 8'hBE;
		16'h2E0: out_word = 8'h28;
		16'h2E1: out_word = 8'h2E;
		16'h2E2: out_word = 8'hEB;
		16'h2E3: out_word = 8'h21;
		16'h2E4: out_word = 8'h04;
		16'h2E5: out_word = 8'h5C;
		16'h2E6: out_word = 8'hBE;
		16'h2E7: out_word = 8'h28;
		16'h2E8: out_word = 8'h27;
		16'h2E9: out_word = 8'hCB;
		16'h2EA: out_word = 8'h7E;
		16'h2EB: out_word = 8'h20;
		16'h2EC: out_word = 8'h04;
		16'h2ED: out_word = 8'hEB;
		16'h2EE: out_word = 8'hCB;
		16'h2EF: out_word = 8'h7E;
		16'h2F0: out_word = 8'hC8;
		16'h2F1: out_word = 8'h5F;
		16'h2F2: out_word = 8'h77;
		16'h2F3: out_word = 8'h23;
		16'h2F4: out_word = 8'h36;
		16'h2F5: out_word = 8'h05;
		16'h2F6: out_word = 8'h23;
		16'h2F7: out_word = 8'h3A;
		16'h2F8: out_word = 8'h09;
		16'h2F9: out_word = 8'h5C;
		16'h2FA: out_word = 8'h77;
		16'h2FB: out_word = 8'h23;
		16'h2FC: out_word = 8'hFD;
		16'h2FD: out_word = 8'h4E;
		16'h2FE: out_word = 8'h07;
		16'h2FF: out_word = 8'hFD;
		16'h300: out_word = 8'h56;
		16'h301: out_word = 8'h01;
		16'h302: out_word = 8'hE5;
		16'h303: out_word = 8'hCD;
		16'h304: out_word = 8'h33;
		16'h305: out_word = 8'h03;
		16'h306: out_word = 8'hE1;
		16'h307: out_word = 8'h77;
		16'h308: out_word = 8'h32;
		16'h309: out_word = 8'h08;
		16'h30A: out_word = 8'h5C;
		16'h30B: out_word = 8'hFD;
		16'h30C: out_word = 8'hCB;
		16'h30D: out_word = 8'h01;
		16'h30E: out_word = 8'hEE;
		16'h30F: out_word = 8'hC9;
		16'h310: out_word = 8'h23;
		16'h311: out_word = 8'h36;
		16'h312: out_word = 8'h05;
		16'h313: out_word = 8'h23;
		16'h314: out_word = 8'h35;
		16'h315: out_word = 8'hC0;
		16'h316: out_word = 8'h3A;
		16'h317: out_word = 8'h0A;
		16'h318: out_word = 8'h5C;
		16'h319: out_word = 8'h77;
		16'h31A: out_word = 8'h23;
		16'h31B: out_word = 8'h7E;
		16'h31C: out_word = 8'h18;
		16'h31D: out_word = 8'hEA;
		16'h31E: out_word = 8'h42;
		16'h31F: out_word = 8'h16;
		16'h320: out_word = 8'h00;
		16'h321: out_word = 8'h7B;
		16'h322: out_word = 8'hFE;
		16'h323: out_word = 8'h27;
		16'h324: out_word = 8'hD0;
		16'h325: out_word = 8'hFE;
		16'h326: out_word = 8'h18;
		16'h327: out_word = 8'h20;
		16'h328: out_word = 8'h03;
		16'h329: out_word = 8'hCB;
		16'h32A: out_word = 8'h78;
		16'h32B: out_word = 8'hC0;
		16'h32C: out_word = 8'h21;
		16'h32D: out_word = 8'h05;
		16'h32E: out_word = 8'h02;
		16'h32F: out_word = 8'h19;
		16'h330: out_word = 8'h7E;
		16'h331: out_word = 8'h37;
		16'h332: out_word = 8'hC9;
		16'h333: out_word = 8'h7B;
		16'h334: out_word = 8'hFE;
		16'h335: out_word = 8'h3A;
		16'h336: out_word = 8'h38;
		16'h337: out_word = 8'h2F;
		16'h338: out_word = 8'h0D;
		16'h339: out_word = 8'hFA;
		16'h33A: out_word = 8'h4F;
		16'h33B: out_word = 8'h03;
		16'h33C: out_word = 8'h28;
		16'h33D: out_word = 8'h03;
		16'h33E: out_word = 8'hC6;
		16'h33F: out_word = 8'h4F;
		16'h340: out_word = 8'hC9;
		16'h341: out_word = 8'h21;
		16'h342: out_word = 8'hEB;
		16'h343: out_word = 8'h01;
		16'h344: out_word = 8'h04;
		16'h345: out_word = 8'h28;
		16'h346: out_word = 8'h03;
		16'h347: out_word = 8'h21;
		16'h348: out_word = 8'h05;
		16'h349: out_word = 8'h02;
		16'h34A: out_word = 8'h16;
		16'h34B: out_word = 8'h00;
		16'h34C: out_word = 8'h19;
		16'h34D: out_word = 8'h7E;
		16'h34E: out_word = 8'hC9;
		16'h34F: out_word = 8'h21;
		16'h350: out_word = 8'h29;
		16'h351: out_word = 8'h02;
		16'h352: out_word = 8'hCB;
		16'h353: out_word = 8'h40;
		16'h354: out_word = 8'h28;
		16'h355: out_word = 8'hF4;
		16'h356: out_word = 8'hCB;
		16'h357: out_word = 8'h5A;
		16'h358: out_word = 8'h28;
		16'h359: out_word = 8'h0A;
		16'h35A: out_word = 8'hFD;
		16'h35B: out_word = 8'hCB;
		16'h35C: out_word = 8'h30;
		16'h35D: out_word = 8'h5E;
		16'h35E: out_word = 8'hC0;
		16'h35F: out_word = 8'h04;
		16'h360: out_word = 8'hC0;
		16'h361: out_word = 8'hC6;
		16'h362: out_word = 8'h20;
		16'h363: out_word = 8'hC9;
		16'h364: out_word = 8'hC6;
		16'h365: out_word = 8'hA5;
		16'h366: out_word = 8'hC9;
		16'h367: out_word = 8'hFE;
		16'h368: out_word = 8'h30;
		16'h369: out_word = 8'hD8;
		16'h36A: out_word = 8'h0D;
		16'h36B: out_word = 8'hFA;
		16'h36C: out_word = 8'h9D;
		16'h36D: out_word = 8'h03;
		16'h36E: out_word = 8'h20;
		16'h36F: out_word = 8'h19;
		16'h370: out_word = 8'h21;
		16'h371: out_word = 8'h54;
		16'h372: out_word = 8'h02;
		16'h373: out_word = 8'hCB;
		16'h374: out_word = 8'h68;
		16'h375: out_word = 8'h28;
		16'h376: out_word = 8'hD3;
		16'h377: out_word = 8'hFE;
		16'h378: out_word = 8'h38;
		16'h379: out_word = 8'h30;
		16'h37A: out_word = 8'h07;
		16'h37B: out_word = 8'hD6;
		16'h37C: out_word = 8'h20;
		16'h37D: out_word = 8'h04;
		16'h37E: out_word = 8'hC8;
		16'h37F: out_word = 8'hC6;
		16'h380: out_word = 8'h08;
		16'h381: out_word = 8'hC9;
		16'h382: out_word = 8'hD6;
		16'h383: out_word = 8'h36;
		16'h384: out_word = 8'h04;
		16'h385: out_word = 8'hC8;
		16'h386: out_word = 8'hC6;
		16'h387: out_word = 8'hFE;
		16'h388: out_word = 8'hC9;
		16'h389: out_word = 8'h21;
		16'h38A: out_word = 8'h30;
		16'h38B: out_word = 8'h02;
		16'h38C: out_word = 8'hFE;
		16'h38D: out_word = 8'h39;
		16'h38E: out_word = 8'h28;
		16'h38F: out_word = 8'hBA;
		16'h390: out_word = 8'hFE;
		16'h391: out_word = 8'h30;
		16'h392: out_word = 8'h28;
		16'h393: out_word = 8'hB6;
		16'h394: out_word = 8'hE6;
		16'h395: out_word = 8'h07;
		16'h396: out_word = 8'hC6;
		16'h397: out_word = 8'h80;
		16'h398: out_word = 8'h04;
		16'h399: out_word = 8'hC8;
		16'h39A: out_word = 8'hEE;
		16'h39B: out_word = 8'h0F;
		16'h39C: out_word = 8'hC9;
		16'h39D: out_word = 8'h04;
		16'h39E: out_word = 8'hC8;
		16'h39F: out_word = 8'hCB;
		16'h3A0: out_word = 8'h68;
		16'h3A1: out_word = 8'h21;
		16'h3A2: out_word = 8'h30;
		16'h3A3: out_word = 8'h02;
		16'h3A4: out_word = 8'h20;
		16'h3A5: out_word = 8'hA4;
		16'h3A6: out_word = 8'hD6;
		16'h3A7: out_word = 8'h10;
		16'h3A8: out_word = 8'hFE;
		16'h3A9: out_word = 8'h22;
		16'h3AA: out_word = 8'h28;
		16'h3AB: out_word = 8'h06;
		16'h3AC: out_word = 8'hFE;
		16'h3AD: out_word = 8'h20;
		16'h3AE: out_word = 8'hC0;
		16'h3AF: out_word = 8'h3E;
		16'h3B0: out_word = 8'h5F;
		16'h3B1: out_word = 8'hC9;
		16'h3B2: out_word = 8'h3E;
		16'h3B3: out_word = 8'h40;
		16'h3B4: out_word = 8'hC9;
		16'h3B5: out_word = 8'hF3;
		16'h3B6: out_word = 8'h7D;
		16'h3B7: out_word = 8'hCB;
		16'h3B8: out_word = 8'h3D;
		16'h3B9: out_word = 8'hCB;
		16'h3BA: out_word = 8'h3D;
		16'h3BB: out_word = 8'h2F;
		16'h3BC: out_word = 8'hE6;
		16'h3BD: out_word = 8'h03;
		16'h3BE: out_word = 8'h4F;
		16'h3BF: out_word = 8'h06;
		16'h3C0: out_word = 8'h00;
		16'h3C1: out_word = 8'hDD;
		16'h3C2: out_word = 8'h21;
		16'h3C3: out_word = 8'hD1;
		16'h3C4: out_word = 8'h03;
		16'h3C5: out_word = 8'hDD;
		16'h3C6: out_word = 8'h09;
		16'h3C7: out_word = 8'h3A;
		16'h3C8: out_word = 8'h48;
		16'h3C9: out_word = 8'h5C;
		16'h3CA: out_word = 8'hE6;
		16'h3CB: out_word = 8'h38;
		16'h3CC: out_word = 8'h0F;
		16'h3CD: out_word = 8'h0F;
		16'h3CE: out_word = 8'h0F;
		16'h3CF: out_word = 8'hF6;
		16'h3D0: out_word = 8'h08;
		16'h3D1: out_word = 8'h00;
		16'h3D2: out_word = 8'h00;
		16'h3D3: out_word = 8'h00;
		16'h3D4: out_word = 8'h04;
		16'h3D5: out_word = 8'h0C;
		16'h3D6: out_word = 8'h0D;
		16'h3D7: out_word = 8'h20;
		16'h3D8: out_word = 8'hFD;
		16'h3D9: out_word = 8'h0E;
		16'h3DA: out_word = 8'h3F;
		16'h3DB: out_word = 8'h05;
		16'h3DC: out_word = 8'hC2;
		16'h3DD: out_word = 8'hD6;
		16'h3DE: out_word = 8'h03;
		16'h3DF: out_word = 8'hEE;
		16'h3E0: out_word = 8'h10;
		16'h3E1: out_word = 8'hD3;
		16'h3E2: out_word = 8'hFE;
		16'h3E3: out_word = 8'h44;
		16'h3E4: out_word = 8'h4F;
		16'h3E5: out_word = 8'hCB;
		16'h3E6: out_word = 8'h67;
		16'h3E7: out_word = 8'h20;
		16'h3E8: out_word = 8'h09;
		16'h3E9: out_word = 8'h7A;
		16'h3EA: out_word = 8'hB3;
		16'h3EB: out_word = 8'h28;
		16'h3EC: out_word = 8'h09;
		16'h3ED: out_word = 8'h79;
		16'h3EE: out_word = 8'h4D;
		16'h3EF: out_word = 8'h1B;
		16'h3F0: out_word = 8'hDD;
		16'h3F1: out_word = 8'hE9;
		16'h3F2: out_word = 8'h4D;
		16'h3F3: out_word = 8'h0C;
		16'h3F4: out_word = 8'hDD;
		16'h3F5: out_word = 8'hE9;
		16'h3F6: out_word = 8'hFB;
		16'h3F7: out_word = 8'hC9;
		16'h3F8: out_word = 8'hEF;
		16'h3F9: out_word = 8'h31;
		16'h3FA: out_word = 8'h27;
		16'h3FB: out_word = 8'hC0;
		16'h3FC: out_word = 8'h03;
		16'h3FD: out_word = 8'h34;
		16'h3FE: out_word = 8'hEC;
		16'h3FF: out_word = 8'h6C;
		16'h400: out_word = 8'h98;
		16'h401: out_word = 8'h1F;
		16'h402: out_word = 8'hF5;
		16'h403: out_word = 8'h04;
		16'h404: out_word = 8'hA1;
		16'h405: out_word = 8'h0F;
		16'h406: out_word = 8'h38;
		16'h407: out_word = 8'h21;
		16'h408: out_word = 8'h92;
		16'h409: out_word = 8'h5C;
		16'h40A: out_word = 8'h7E;
		16'h40B: out_word = 8'hA7;
		16'h40C: out_word = 8'h20;
		16'h40D: out_word = 8'h5E;
		16'h40E: out_word = 8'h23;
		16'h40F: out_word = 8'h4E;
		16'h410: out_word = 8'h23;
		16'h411: out_word = 8'h46;
		16'h412: out_word = 8'h78;
		16'h413: out_word = 8'h17;
		16'h414: out_word = 8'h9F;
		16'h415: out_word = 8'hB9;
		16'h416: out_word = 8'h20;
		16'h417: out_word = 8'h54;
		16'h418: out_word = 8'h23;
		16'h419: out_word = 8'hBE;
		16'h41A: out_word = 8'h20;
		16'h41B: out_word = 8'h50;
		16'h41C: out_word = 8'h78;
		16'h41D: out_word = 8'hC6;
		16'h41E: out_word = 8'h3C;
		16'h41F: out_word = 8'hF2;
		16'h420: out_word = 8'h25;
		16'h421: out_word = 8'h04;
		16'h422: out_word = 8'hE2;
		16'h423: out_word = 8'h6C;
		16'h424: out_word = 8'h04;
		16'h425: out_word = 8'h06;
		16'h426: out_word = 8'hFA;
		16'h427: out_word = 8'h04;
		16'h428: out_word = 8'hD6;
		16'h429: out_word = 8'h0C;
		16'h42A: out_word = 8'h30;
		16'h42B: out_word = 8'hFB;
		16'h42C: out_word = 8'hC6;
		16'h42D: out_word = 8'h0C;
		16'h42E: out_word = 8'hC5;
		16'h42F: out_word = 8'h21;
		16'h430: out_word = 8'h6E;
		16'h431: out_word = 8'h04;
		16'h432: out_word = 8'hCD;
		16'h433: out_word = 8'h06;
		16'h434: out_word = 8'h34;
		16'h435: out_word = 8'hCD;
		16'h436: out_word = 8'hB4;
		16'h437: out_word = 8'h33;
		16'h438: out_word = 8'hEF;
		16'h439: out_word = 8'h04;
		16'h43A: out_word = 8'h38;
		16'h43B: out_word = 8'hF1;
		16'h43C: out_word = 8'h86;
		16'h43D: out_word = 8'h77;
		16'h43E: out_word = 8'hEF;
		16'h43F: out_word = 8'hC0;
		16'h440: out_word = 8'h02;
		16'h441: out_word = 8'h31;
		16'h442: out_word = 8'h38;
		16'h443: out_word = 8'hCD;
		16'h444: out_word = 8'h94;
		16'h445: out_word = 8'h1E;
		16'h446: out_word = 8'hFE;
		16'h447: out_word = 8'h0B;
		16'h448: out_word = 8'h30;
		16'h449: out_word = 8'h22;
		16'h44A: out_word = 8'hEF;
		16'h44B: out_word = 8'hE0;
		16'h44C: out_word = 8'h04;
		16'h44D: out_word = 8'hE0;
		16'h44E: out_word = 8'h34;
		16'h44F: out_word = 8'h80;
		16'h450: out_word = 8'h43;
		16'h451: out_word = 8'h55;
		16'h452: out_word = 8'h9F;
		16'h453: out_word = 8'h80;
		16'h454: out_word = 8'h01;
		16'h455: out_word = 8'h05;
		16'h456: out_word = 8'h34;
		16'h457: out_word = 8'h35;
		16'h458: out_word = 8'h71;
		16'h459: out_word = 8'h03;
		16'h45A: out_word = 8'h38;
		16'h45B: out_word = 8'hCD;
		16'h45C: out_word = 8'h99;
		16'h45D: out_word = 8'h1E;
		16'h45E: out_word = 8'hC5;
		16'h45F: out_word = 8'hCD;
		16'h460: out_word = 8'h99;
		16'h461: out_word = 8'h1E;
		16'h462: out_word = 8'hE1;
		16'h463: out_word = 8'h50;
		16'h464: out_word = 8'h59;
		16'h465: out_word = 8'h7A;
		16'h466: out_word = 8'hB3;
		16'h467: out_word = 8'hC8;
		16'h468: out_word = 8'h1B;
		16'h469: out_word = 8'hC3;
		16'h46A: out_word = 8'hB5;
		16'h46B: out_word = 8'h03;
		16'h46C: out_word = 8'hCF;
		16'h46D: out_word = 8'h0A;
		16'h46E: out_word = 8'h89;
		16'h46F: out_word = 8'h02;
		16'h470: out_word = 8'hD0;
		16'h471: out_word = 8'h12;
		16'h472: out_word = 8'h86;
		16'h473: out_word = 8'h89;
		16'h474: out_word = 8'h0A;
		16'h475: out_word = 8'h97;
		16'h476: out_word = 8'h60;
		16'h477: out_word = 8'h75;
		16'h478: out_word = 8'h89;
		16'h479: out_word = 8'h12;
		16'h47A: out_word = 8'hD5;
		16'h47B: out_word = 8'h17;
		16'h47C: out_word = 8'h1F;
		16'h47D: out_word = 8'h89;
		16'h47E: out_word = 8'h1B;
		16'h47F: out_word = 8'h90;
		16'h480: out_word = 8'h41;
		16'h481: out_word = 8'h02;
		16'h482: out_word = 8'h89;
		16'h483: out_word = 8'h24;
		16'h484: out_word = 8'hD0;
		16'h485: out_word = 8'h53;
		16'h486: out_word = 8'hCA;
		16'h487: out_word = 8'h89;
		16'h488: out_word = 8'h2E;
		16'h489: out_word = 8'h9D;
		16'h48A: out_word = 8'h36;
		16'h48B: out_word = 8'hB1;
		16'h48C: out_word = 8'h89;
		16'h48D: out_word = 8'h38;
		16'h48E: out_word = 8'hFF;
		16'h48F: out_word = 8'h49;
		16'h490: out_word = 8'h3E;
		16'h491: out_word = 8'h89;
		16'h492: out_word = 8'h43;
		16'h493: out_word = 8'hFF;
		16'h494: out_word = 8'h6A;
		16'h495: out_word = 8'h73;
		16'h496: out_word = 8'h89;
		16'h497: out_word = 8'h4F;
		16'h498: out_word = 8'hA7;
		16'h499: out_word = 8'h00;
		16'h49A: out_word = 8'h54;
		16'h49B: out_word = 8'h89;
		16'h49C: out_word = 8'h5C;
		16'h49D: out_word = 8'h00;
		16'h49E: out_word = 8'h00;
		16'h49F: out_word = 8'h00;
		16'h4A0: out_word = 8'h89;
		16'h4A1: out_word = 8'h69;
		16'h4A2: out_word = 8'h14;
		16'h4A3: out_word = 8'hF6;
		16'h4A4: out_word = 8'h24;
		16'h4A5: out_word = 8'h89;
		16'h4A6: out_word = 8'h76;
		16'h4A7: out_word = 8'hF1;
		16'h4A8: out_word = 8'h10;
		16'h4A9: out_word = 8'h05;
		16'h4AA: out_word = 8'hCD;
		16'h4AB: out_word = 8'hFB;
		16'h4AC: out_word = 8'h24;
		16'h4AD: out_word = 8'h3A;
		16'h4AE: out_word = 8'h3B;
		16'h4AF: out_word = 8'h5C;
		16'h4B0: out_word = 8'h87;
		16'h4B1: out_word = 8'hFA;
		16'h4B2: out_word = 8'h8A;
		16'h4B3: out_word = 8'h1C;
		16'h4B4: out_word = 8'hE1;
		16'h4B5: out_word = 8'hD0;
		16'h4B6: out_word = 8'hE5;
		16'h4B7: out_word = 8'hCD;
		16'h4B8: out_word = 8'hF1;
		16'h4B9: out_word = 8'h2B;
		16'h4BA: out_word = 8'h62;
		16'h4BB: out_word = 8'h6B;
		16'h4BC: out_word = 8'h0D;
		16'h4BD: out_word = 8'hF8;
		16'h4BE: out_word = 8'h09;
		16'h4BF: out_word = 8'hCB;
		16'h4C0: out_word = 8'hFE;
		16'h4C1: out_word = 8'hC9;
		16'h4C2: out_word = 8'h21;
		16'h4C3: out_word = 8'h3F;
		16'h4C4: out_word = 8'h05;
		16'h4C5: out_word = 8'hE5;
		16'h4C6: out_word = 8'h21;
		16'h4C7: out_word = 8'h80;
		16'h4C8: out_word = 8'h1F;
		16'h4C9: out_word = 8'hCB;
		16'h4CA: out_word = 8'h7F;
		16'h4CB: out_word = 8'h28;
		16'h4CC: out_word = 8'h03;
		16'h4CD: out_word = 8'h21;
		16'h4CE: out_word = 8'h98;
		16'h4CF: out_word = 8'h0C;
		16'h4D0: out_word = 8'h08;
		16'h4D1: out_word = 8'h13;
		16'h4D2: out_word = 8'hDD;
		16'h4D3: out_word = 8'h2B;
		16'h4D4: out_word = 8'hF3;
		16'h4D5: out_word = 8'h3E;
		16'h4D6: out_word = 8'h02;
		16'h4D7: out_word = 8'h47;
		16'h4D8: out_word = 8'h10;
		16'h4D9: out_word = 8'hFE;
		16'h4DA: out_word = 8'hD3;
		16'h4DB: out_word = 8'hFE;
		16'h4DC: out_word = 8'hEE;
		16'h4DD: out_word = 8'h0F;
		16'h4DE: out_word = 8'h06;
		16'h4DF: out_word = 8'hA4;
		16'h4E0: out_word = 8'h2D;
		16'h4E1: out_word = 8'h20;
		16'h4E2: out_word = 8'hF5;
		16'h4E3: out_word = 8'h05;
		16'h4E4: out_word = 8'h25;
		16'h4E5: out_word = 8'hF2;
		16'h4E6: out_word = 8'hD8;
		16'h4E7: out_word = 8'h04;
		16'h4E8: out_word = 8'h06;
		16'h4E9: out_word = 8'h2F;
		16'h4EA: out_word = 8'h10;
		16'h4EB: out_word = 8'hFE;
		16'h4EC: out_word = 8'hD3;
		16'h4ED: out_word = 8'hFE;
		16'h4EE: out_word = 8'h3E;
		16'h4EF: out_word = 8'h0D;
		16'h4F0: out_word = 8'h06;
		16'h4F1: out_word = 8'h37;
		16'h4F2: out_word = 8'h10;
		16'h4F3: out_word = 8'hFE;
		16'h4F4: out_word = 8'hD3;
		16'h4F5: out_word = 8'hFE;
		16'h4F6: out_word = 8'h01;
		16'h4F7: out_word = 8'h0E;
		16'h4F8: out_word = 8'h3B;
		16'h4F9: out_word = 8'h08;
		16'h4FA: out_word = 8'h6F;
		16'h4FB: out_word = 8'hC3;
		16'h4FC: out_word = 8'h07;
		16'h4FD: out_word = 8'h05;
		16'h4FE: out_word = 8'h7A;
		16'h4FF: out_word = 8'hB3;
		16'h500: out_word = 8'h28;
		16'h501: out_word = 8'h0C;
		16'h502: out_word = 8'hDD;
		16'h503: out_word = 8'h6E;
		16'h504: out_word = 8'h00;
		16'h505: out_word = 8'h7C;
		16'h506: out_word = 8'hAD;
		16'h507: out_word = 8'h67;
		16'h508: out_word = 8'h3E;
		16'h509: out_word = 8'h01;
		16'h50A: out_word = 8'h37;
		16'h50B: out_word = 8'hC3;
		16'h50C: out_word = 8'h25;
		16'h50D: out_word = 8'h05;
		16'h50E: out_word = 8'h6C;
		16'h50F: out_word = 8'h18;
		16'h510: out_word = 8'hF4;
		16'h511: out_word = 8'h79;
		16'h512: out_word = 8'hCB;
		16'h513: out_word = 8'h78;
		16'h514: out_word = 8'h10;
		16'h515: out_word = 8'hFE;
		16'h516: out_word = 8'h30;
		16'h517: out_word = 8'h04;
		16'h518: out_word = 8'h06;
		16'h519: out_word = 8'h42;
		16'h51A: out_word = 8'h10;
		16'h51B: out_word = 8'hFE;
		16'h51C: out_word = 8'hD3;
		16'h51D: out_word = 8'hFE;
		16'h51E: out_word = 8'h06;
		16'h51F: out_word = 8'h3E;
		16'h520: out_word = 8'h20;
		16'h521: out_word = 8'hEF;
		16'h522: out_word = 8'h05;
		16'h523: out_word = 8'hAF;
		16'h524: out_word = 8'h3C;
		16'h525: out_word = 8'hCB;
		16'h526: out_word = 8'h15;
		16'h527: out_word = 8'hC2;
		16'h528: out_word = 8'h14;
		16'h529: out_word = 8'h05;
		16'h52A: out_word = 8'h1B;
		16'h52B: out_word = 8'hDD;
		16'h52C: out_word = 8'h23;
		16'h52D: out_word = 8'h06;
		16'h52E: out_word = 8'h31;
		16'h52F: out_word = 8'h3E;
		16'h530: out_word = 8'h7F;
		16'h531: out_word = 8'hDB;
		16'h532: out_word = 8'hFE;
		16'h533: out_word = 8'h1F;
		16'h534: out_word = 8'hD0;
		16'h535: out_word = 8'h7A;
		16'h536: out_word = 8'h3C;
		16'h537: out_word = 8'hC2;
		16'h538: out_word = 8'hFE;
		16'h539: out_word = 8'h04;
		16'h53A: out_word = 8'h06;
		16'h53B: out_word = 8'h3B;
		16'h53C: out_word = 8'h10;
		16'h53D: out_word = 8'hFE;
		16'h53E: out_word = 8'hC9;
		16'h53F: out_word = 8'hF5;
		16'h540: out_word = 8'h3A;
		16'h541: out_word = 8'h48;
		16'h542: out_word = 8'h5C;
		16'h543: out_word = 8'hE6;
		16'h544: out_word = 8'h38;
		16'h545: out_word = 8'h0F;
		16'h546: out_word = 8'h0F;
		16'h547: out_word = 8'h0F;
		16'h548: out_word = 8'hD3;
		16'h549: out_word = 8'hFE;
		16'h54A: out_word = 8'h3E;
		16'h54B: out_word = 8'h7F;
		16'h54C: out_word = 8'hDB;
		16'h54D: out_word = 8'hFE;
		16'h54E: out_word = 8'h1F;
		16'h54F: out_word = 8'hFB;
		16'h550: out_word = 8'h38;
		16'h551: out_word = 8'h02;
		16'h552: out_word = 8'hCF;
		16'h553: out_word = 8'h0C;
		16'h554: out_word = 8'hF1;
		16'h555: out_word = 8'hC9;
		16'h556: out_word = 8'h14;
		16'h557: out_word = 8'h08;
		16'h558: out_word = 8'h15;
		16'h559: out_word = 8'hF3;
		16'h55A: out_word = 8'h3E;
		16'h55B: out_word = 8'h0F;
		16'h55C: out_word = 8'hD3;
		16'h55D: out_word = 8'hFE;
		16'h55E: out_word = 8'h21;
		16'h55F: out_word = 8'h3F;
		16'h560: out_word = 8'h05;
		16'h561: out_word = 8'hE5;
		16'h562: out_word = 8'hDB;
		16'h563: out_word = 8'hFE;
		16'h564: out_word = 8'h1F;
		16'h565: out_word = 8'hE6;
		16'h566: out_word = 8'h20;
		16'h567: out_word = 8'hF6;
		16'h568: out_word = 8'h02;
		16'h569: out_word = 8'h4F;
		16'h56A: out_word = 8'hBF;
		16'h56B: out_word = 8'hC0;
		16'h56C: out_word = 8'hCD;
		16'h56D: out_word = 8'hE7;
		16'h56E: out_word = 8'h05;
		16'h56F: out_word = 8'h30;
		16'h570: out_word = 8'hFA;
		16'h571: out_word = 8'h21;
		16'h572: out_word = 8'h15;
		16'h573: out_word = 8'h04;
		16'h574: out_word = 8'h10;
		16'h575: out_word = 8'hFE;
		16'h576: out_word = 8'h2B;
		16'h577: out_word = 8'h7C;
		16'h578: out_word = 8'hB5;
		16'h579: out_word = 8'h20;
		16'h57A: out_word = 8'hF9;
		16'h57B: out_word = 8'hCD;
		16'h57C: out_word = 8'hE3;
		16'h57D: out_word = 8'h05;
		16'h57E: out_word = 8'h30;
		16'h57F: out_word = 8'hEB;
		16'h580: out_word = 8'h06;
		16'h581: out_word = 8'h9C;
		16'h582: out_word = 8'hCD;
		16'h583: out_word = 8'hE3;
		16'h584: out_word = 8'h05;
		16'h585: out_word = 8'h30;
		16'h586: out_word = 8'hE4;
		16'h587: out_word = 8'h3E;
		16'h588: out_word = 8'hC6;
		16'h589: out_word = 8'hB8;
		16'h58A: out_word = 8'h30;
		16'h58B: out_word = 8'hE0;
		16'h58C: out_word = 8'h24;
		16'h58D: out_word = 8'h20;
		16'h58E: out_word = 8'hF1;
		16'h58F: out_word = 8'h06;
		16'h590: out_word = 8'hC9;
		16'h591: out_word = 8'hCD;
		16'h592: out_word = 8'hE7;
		16'h593: out_word = 8'h05;
		16'h594: out_word = 8'h30;
		16'h595: out_word = 8'hD5;
		16'h596: out_word = 8'h78;
		16'h597: out_word = 8'hFE;
		16'h598: out_word = 8'hD4;
		16'h599: out_word = 8'h30;
		16'h59A: out_word = 8'hF4;
		16'h59B: out_word = 8'hCD;
		16'h59C: out_word = 8'hE7;
		16'h59D: out_word = 8'h05;
		16'h59E: out_word = 8'hD0;
		16'h59F: out_word = 8'h79;
		16'h5A0: out_word = 8'hEE;
		16'h5A1: out_word = 8'h03;
		16'h5A2: out_word = 8'h4F;
		16'h5A3: out_word = 8'h26;
		16'h5A4: out_word = 8'h00;
		16'h5A5: out_word = 8'h06;
		16'h5A6: out_word = 8'hB0;
		16'h5A7: out_word = 8'h18;
		16'h5A8: out_word = 8'h1F;
		16'h5A9: out_word = 8'h08;
		16'h5AA: out_word = 8'h20;
		16'h5AB: out_word = 8'h07;
		16'h5AC: out_word = 8'h30;
		16'h5AD: out_word = 8'h0F;
		16'h5AE: out_word = 8'hDD;
		16'h5AF: out_word = 8'h75;
		16'h5B0: out_word = 8'h00;
		16'h5B1: out_word = 8'h18;
		16'h5B2: out_word = 8'h0F;
		16'h5B3: out_word = 8'hCB;
		16'h5B4: out_word = 8'h11;
		16'h5B5: out_word = 8'hAD;
		16'h5B6: out_word = 8'hC0;
		16'h5B7: out_word = 8'h79;
		16'h5B8: out_word = 8'h1F;
		16'h5B9: out_word = 8'h4F;
		16'h5BA: out_word = 8'h13;
		16'h5BB: out_word = 8'h18;
		16'h5BC: out_word = 8'h07;
		16'h5BD: out_word = 8'hDD;
		16'h5BE: out_word = 8'h7E;
		16'h5BF: out_word = 8'h00;
		16'h5C0: out_word = 8'hAD;
		16'h5C1: out_word = 8'hC0;
		16'h5C2: out_word = 8'hDD;
		16'h5C3: out_word = 8'h23;
		16'h5C4: out_word = 8'h1B;
		16'h5C5: out_word = 8'h08;
		16'h5C6: out_word = 8'h06;
		16'h5C7: out_word = 8'hB2;
		16'h5C8: out_word = 8'h2E;
		16'h5C9: out_word = 8'h01;
		16'h5CA: out_word = 8'hCD;
		16'h5CB: out_word = 8'hE3;
		16'h5CC: out_word = 8'h05;
		16'h5CD: out_word = 8'hD0;
		16'h5CE: out_word = 8'h3E;
		16'h5CF: out_word = 8'hCB;
		16'h5D0: out_word = 8'hB8;
		16'h5D1: out_word = 8'hCB;
		16'h5D2: out_word = 8'h15;
		16'h5D3: out_word = 8'h06;
		16'h5D4: out_word = 8'hB0;
		16'h5D5: out_word = 8'hD2;
		16'h5D6: out_word = 8'hCA;
		16'h5D7: out_word = 8'h05;
		16'h5D8: out_word = 8'h7C;
		16'h5D9: out_word = 8'hAD;
		16'h5DA: out_word = 8'h67;
		16'h5DB: out_word = 8'h7A;
		16'h5DC: out_word = 8'hB3;
		16'h5DD: out_word = 8'h20;
		16'h5DE: out_word = 8'hCA;
		16'h5DF: out_word = 8'h7C;
		16'h5E0: out_word = 8'hFE;
		16'h5E1: out_word = 8'h01;
		16'h5E2: out_word = 8'hC9;
		16'h5E3: out_word = 8'hCD;
		16'h5E4: out_word = 8'hE7;
		16'h5E5: out_word = 8'h05;
		16'h5E6: out_word = 8'hD0;
		16'h5E7: out_word = 8'h3E;
		16'h5E8: out_word = 8'h16;
		16'h5E9: out_word = 8'h3D;
		16'h5EA: out_word = 8'h20;
		16'h5EB: out_word = 8'hFD;
		16'h5EC: out_word = 8'hA7;
		16'h5ED: out_word = 8'h04;
		16'h5EE: out_word = 8'hC8;
		16'h5EF: out_word = 8'h3E;
		16'h5F0: out_word = 8'h7F;
		16'h5F1: out_word = 8'hDB;
		16'h5F2: out_word = 8'hFE;
		16'h5F3: out_word = 8'h1F;
		16'h5F4: out_word = 8'hD0;
		16'h5F5: out_word = 8'hA9;
		16'h5F6: out_word = 8'hE6;
		16'h5F7: out_word = 8'h20;
		16'h5F8: out_word = 8'h28;
		16'h5F9: out_word = 8'hF3;
		16'h5FA: out_word = 8'h79;
		16'h5FB: out_word = 8'h2F;
		16'h5FC: out_word = 8'h4F;
		16'h5FD: out_word = 8'hE6;
		16'h5FE: out_word = 8'h07;
		16'h5FF: out_word = 8'hF6;
		16'h600: out_word = 8'h08;
		16'h601: out_word = 8'hD3;
		16'h602: out_word = 8'hFE;
		16'h603: out_word = 8'h37;
		16'h604: out_word = 8'hC9;
		16'h605: out_word = 8'hF1;
		16'h606: out_word = 8'h3A;
		16'h607: out_word = 8'h74;
		16'h608: out_word = 8'h5C;
		16'h609: out_word = 8'hD6;
		16'h60A: out_word = 8'hE0;
		16'h60B: out_word = 8'h32;
		16'h60C: out_word = 8'h74;
		16'h60D: out_word = 8'h5C;
		16'h60E: out_word = 8'hCD;
		16'h60F: out_word = 8'h8C;
		16'h610: out_word = 8'h1C;
		16'h611: out_word = 8'hCD;
		16'h612: out_word = 8'h30;
		16'h613: out_word = 8'h25;
		16'h614: out_word = 8'h28;
		16'h615: out_word = 8'h3C;
		16'h616: out_word = 8'h01;
		16'h617: out_word = 8'h11;
		16'h618: out_word = 8'h00;
		16'h619: out_word = 8'h3A;
		16'h61A: out_word = 8'h74;
		16'h61B: out_word = 8'h5C;
		16'h61C: out_word = 8'hA7;
		16'h61D: out_word = 8'h28;
		16'h61E: out_word = 8'h02;
		16'h61F: out_word = 8'h0E;
		16'h620: out_word = 8'h22;
		16'h621: out_word = 8'hF7;
		16'h622: out_word = 8'hD5;
		16'h623: out_word = 8'hDD;
		16'h624: out_word = 8'hE1;
		16'h625: out_word = 8'h06;
		16'h626: out_word = 8'h0B;
		16'h627: out_word = 8'h3E;
		16'h628: out_word = 8'h20;
		16'h629: out_word = 8'h12;
		16'h62A: out_word = 8'h13;
		16'h62B: out_word = 8'h10;
		16'h62C: out_word = 8'hFC;
		16'h62D: out_word = 8'hDD;
		16'h62E: out_word = 8'h36;
		16'h62F: out_word = 8'h01;
		16'h630: out_word = 8'hFF;
		16'h631: out_word = 8'hCD;
		16'h632: out_word = 8'hF1;
		16'h633: out_word = 8'h2B;
		16'h634: out_word = 8'h21;
		16'h635: out_word = 8'hF6;
		16'h636: out_word = 8'hFF;
		16'h637: out_word = 8'h0B;
		16'h638: out_word = 8'h09;
		16'h639: out_word = 8'h03;
		16'h63A: out_word = 8'h30;
		16'h63B: out_word = 8'h0F;
		16'h63C: out_word = 8'h3A;
		16'h63D: out_word = 8'h74;
		16'h63E: out_word = 8'h5C;
		16'h63F: out_word = 8'hA7;
		16'h640: out_word = 8'h20;
		16'h641: out_word = 8'h02;
		16'h642: out_word = 8'hCF;
		16'h643: out_word = 8'h0E;
		16'h644: out_word = 8'h78;
		16'h645: out_word = 8'hB1;
		16'h646: out_word = 8'h28;
		16'h647: out_word = 8'h0A;
		16'h648: out_word = 8'h01;
		16'h649: out_word = 8'h0A;
		16'h64A: out_word = 8'h00;
		16'h64B: out_word = 8'hDD;
		16'h64C: out_word = 8'hE5;
		16'h64D: out_word = 8'hE1;
		16'h64E: out_word = 8'h23;
		16'h64F: out_word = 8'hEB;
		16'h650: out_word = 8'hED;
		16'h651: out_word = 8'hB0;
		16'h652: out_word = 8'hDF;
		16'h653: out_word = 8'hFE;
		16'h654: out_word = 8'hE4;
		16'h655: out_word = 8'h20;
		16'h656: out_word = 8'h49;
		16'h657: out_word = 8'h3A;
		16'h658: out_word = 8'h74;
		16'h659: out_word = 8'h5C;
		16'h65A: out_word = 8'hFE;
		16'h65B: out_word = 8'h03;
		16'h65C: out_word = 8'hCA;
		16'h65D: out_word = 8'h8A;
		16'h65E: out_word = 8'h1C;
		16'h65F: out_word = 8'hE7;
		16'h660: out_word = 8'hCD;
		16'h661: out_word = 8'hB2;
		16'h662: out_word = 8'h28;
		16'h663: out_word = 8'hCB;
		16'h664: out_word = 8'hF9;
		16'h665: out_word = 8'h30;
		16'h666: out_word = 8'h0B;
		16'h667: out_word = 8'h21;
		16'h668: out_word = 8'h00;
		16'h669: out_word = 8'h00;
		16'h66A: out_word = 8'h3A;
		16'h66B: out_word = 8'h74;
		16'h66C: out_word = 8'h5C;
		16'h66D: out_word = 8'h3D;
		16'h66E: out_word = 8'h28;
		16'h66F: out_word = 8'h15;
		16'h670: out_word = 8'hCF;
		16'h671: out_word = 8'h01;
		16'h672: out_word = 8'hC2;
		16'h673: out_word = 8'h8A;
		16'h674: out_word = 8'h1C;
		16'h675: out_word = 8'hCD;
		16'h676: out_word = 8'h30;
		16'h677: out_word = 8'h25;
		16'h678: out_word = 8'h28;
		16'h679: out_word = 8'h18;
		16'h67A: out_word = 8'h23;
		16'h67B: out_word = 8'h7E;
		16'h67C: out_word = 8'hDD;
		16'h67D: out_word = 8'h77;
		16'h67E: out_word = 8'h0B;
		16'h67F: out_word = 8'h23;
		16'h680: out_word = 8'h7E;
		16'h681: out_word = 8'hDD;
		16'h682: out_word = 8'h77;
		16'h683: out_word = 8'h0C;
		16'h684: out_word = 8'h23;
		16'h685: out_word = 8'hDD;
		16'h686: out_word = 8'h71;
		16'h687: out_word = 8'h0E;
		16'h688: out_word = 8'h3E;
		16'h689: out_word = 8'h01;
		16'h68A: out_word = 8'hCB;
		16'h68B: out_word = 8'h71;
		16'h68C: out_word = 8'h28;
		16'h68D: out_word = 8'h01;
		16'h68E: out_word = 8'h3C;
		16'h68F: out_word = 8'hDD;
		16'h690: out_word = 8'h77;
		16'h691: out_word = 8'h00;
		16'h692: out_word = 8'hEB;
		16'h693: out_word = 8'hE7;
		16'h694: out_word = 8'hFE;
		16'h695: out_word = 8'h29;
		16'h696: out_word = 8'h20;
		16'h697: out_word = 8'hDA;
		16'h698: out_word = 8'hE7;
		16'h699: out_word = 8'hCD;
		16'h69A: out_word = 8'hEE;
		16'h69B: out_word = 8'h1B;
		16'h69C: out_word = 8'hEB;
		16'h69D: out_word = 8'hC3;
		16'h69E: out_word = 8'h5A;
		16'h69F: out_word = 8'h07;
		16'h6A0: out_word = 8'hFE;
		16'h6A1: out_word = 8'hAA;
		16'h6A2: out_word = 8'h20;
		16'h6A3: out_word = 8'h1F;
		16'h6A4: out_word = 8'h3A;
		16'h6A5: out_word = 8'h74;
		16'h6A6: out_word = 8'h5C;
		16'h6A7: out_word = 8'hFE;
		16'h6A8: out_word = 8'h03;
		16'h6A9: out_word = 8'hCA;
		16'h6AA: out_word = 8'h8A;
		16'h6AB: out_word = 8'h1C;
		16'h6AC: out_word = 8'hE7;
		16'h6AD: out_word = 8'hCD;
		16'h6AE: out_word = 8'hEE;
		16'h6AF: out_word = 8'h1B;
		16'h6B0: out_word = 8'hDD;
		16'h6B1: out_word = 8'h36;
		16'h6B2: out_word = 8'h0B;
		16'h6B3: out_word = 8'h00;
		16'h6B4: out_word = 8'hDD;
		16'h6B5: out_word = 8'h36;
		16'h6B6: out_word = 8'h0C;
		16'h6B7: out_word = 8'h1B;
		16'h6B8: out_word = 8'h21;
		16'h6B9: out_word = 8'h00;
		16'h6BA: out_word = 8'h40;
		16'h6BB: out_word = 8'hDD;
		16'h6BC: out_word = 8'h75;
		16'h6BD: out_word = 8'h0D;
		16'h6BE: out_word = 8'hDD;
		16'h6BF: out_word = 8'h74;
		16'h6C0: out_word = 8'h0E;
		16'h6C1: out_word = 8'h18;
		16'h6C2: out_word = 8'h4D;
		16'h6C3: out_word = 8'hFE;
		16'h6C4: out_word = 8'hAF;
		16'h6C5: out_word = 8'h20;
		16'h6C6: out_word = 8'h4F;
		16'h6C7: out_word = 8'h3A;
		16'h6C8: out_word = 8'h74;
		16'h6C9: out_word = 8'h5C;
		16'h6CA: out_word = 8'hFE;
		16'h6CB: out_word = 8'h03;
		16'h6CC: out_word = 8'hCA;
		16'h6CD: out_word = 8'h8A;
		16'h6CE: out_word = 8'h1C;
		16'h6CF: out_word = 8'hE7;
		16'h6D0: out_word = 8'hCD;
		16'h6D1: out_word = 8'h48;
		16'h6D2: out_word = 8'h20;
		16'h6D3: out_word = 8'h20;
		16'h6D4: out_word = 8'h0C;
		16'h6D5: out_word = 8'h3A;
		16'h6D6: out_word = 8'h74;
		16'h6D7: out_word = 8'h5C;
		16'h6D8: out_word = 8'hA7;
		16'h6D9: out_word = 8'hCA;
		16'h6DA: out_word = 8'h8A;
		16'h6DB: out_word = 8'h1C;
		16'h6DC: out_word = 8'hCD;
		16'h6DD: out_word = 8'hE6;
		16'h6DE: out_word = 8'h1C;
		16'h6DF: out_word = 8'h18;
		16'h6E0: out_word = 8'h0F;
		16'h6E1: out_word = 8'hCD;
		16'h6E2: out_word = 8'h82;
		16'h6E3: out_word = 8'h1C;
		16'h6E4: out_word = 8'hDF;
		16'h6E5: out_word = 8'hFE;
		16'h6E6: out_word = 8'h2C;
		16'h6E7: out_word = 8'h28;
		16'h6E8: out_word = 8'h0C;
		16'h6E9: out_word = 8'h3A;
		16'h6EA: out_word = 8'h74;
		16'h6EB: out_word = 8'h5C;
		16'h6EC: out_word = 8'hA7;
		16'h6ED: out_word = 8'hCA;
		16'h6EE: out_word = 8'h8A;
		16'h6EF: out_word = 8'h1C;
		16'h6F0: out_word = 8'hCD;
		16'h6F1: out_word = 8'hE6;
		16'h6F2: out_word = 8'h1C;
		16'h6F3: out_word = 8'h18;
		16'h6F4: out_word = 8'h04;
		16'h6F5: out_word = 8'hE7;
		16'h6F6: out_word = 8'hCD;
		16'h6F7: out_word = 8'h82;
		16'h6F8: out_word = 8'h1C;
		16'h6F9: out_word = 8'hCD;
		16'h6FA: out_word = 8'hEE;
		16'h6FB: out_word = 8'h1B;
		16'h6FC: out_word = 8'hCD;
		16'h6FD: out_word = 8'h99;
		16'h6FE: out_word = 8'h1E;
		16'h6FF: out_word = 8'hDD;
		16'h700: out_word = 8'h71;
		16'h701: out_word = 8'h0B;
		16'h702: out_word = 8'hDD;
		16'h703: out_word = 8'h70;
		16'h704: out_word = 8'h0C;
		16'h705: out_word = 8'hCD;
		16'h706: out_word = 8'h99;
		16'h707: out_word = 8'h1E;
		16'h708: out_word = 8'hDD;
		16'h709: out_word = 8'h71;
		16'h70A: out_word = 8'h0D;
		16'h70B: out_word = 8'hDD;
		16'h70C: out_word = 8'h70;
		16'h70D: out_word = 8'h0E;
		16'h70E: out_word = 8'h60;
		16'h70F: out_word = 8'h69;
		16'h710: out_word = 8'hDD;
		16'h711: out_word = 8'h36;
		16'h712: out_word = 8'h00;
		16'h713: out_word = 8'h03;
		16'h714: out_word = 8'h18;
		16'h715: out_word = 8'h44;
		16'h716: out_word = 8'hFE;
		16'h717: out_word = 8'hCA;
		16'h718: out_word = 8'h28;
		16'h719: out_word = 8'h09;
		16'h71A: out_word = 8'hCD;
		16'h71B: out_word = 8'hEE;
		16'h71C: out_word = 8'h1B;
		16'h71D: out_word = 8'hDD;
		16'h71E: out_word = 8'h36;
		16'h71F: out_word = 8'h0E;
		16'h720: out_word = 8'h80;
		16'h721: out_word = 8'h18;
		16'h722: out_word = 8'h17;
		16'h723: out_word = 8'h3A;
		16'h724: out_word = 8'h74;
		16'h725: out_word = 8'h5C;
		16'h726: out_word = 8'hA7;
		16'h727: out_word = 8'hC2;
		16'h728: out_word = 8'h8A;
		16'h729: out_word = 8'h1C;
		16'h72A: out_word = 8'hE7;
		16'h72B: out_word = 8'hCD;
		16'h72C: out_word = 8'h82;
		16'h72D: out_word = 8'h1C;
		16'h72E: out_word = 8'hCD;
		16'h72F: out_word = 8'hEE;
		16'h730: out_word = 8'h1B;
		16'h731: out_word = 8'hCD;
		16'h732: out_word = 8'h99;
		16'h733: out_word = 8'h1E;
		16'h734: out_word = 8'hDD;
		16'h735: out_word = 8'h71;
		16'h736: out_word = 8'h0D;
		16'h737: out_word = 8'hDD;
		16'h738: out_word = 8'h70;
		16'h739: out_word = 8'h0E;
		16'h73A: out_word = 8'hDD;
		16'h73B: out_word = 8'h36;
		16'h73C: out_word = 8'h00;
		16'h73D: out_word = 8'h00;
		16'h73E: out_word = 8'h2A;
		16'h73F: out_word = 8'h59;
		16'h740: out_word = 8'h5C;
		16'h741: out_word = 8'hED;
		16'h742: out_word = 8'h5B;
		16'h743: out_word = 8'h53;
		16'h744: out_word = 8'h5C;
		16'h745: out_word = 8'h37;
		16'h746: out_word = 8'hED;
		16'h747: out_word = 8'h52;
		16'h748: out_word = 8'hDD;
		16'h749: out_word = 8'h75;
		16'h74A: out_word = 8'h0B;
		16'h74B: out_word = 8'hDD;
		16'h74C: out_word = 8'h74;
		16'h74D: out_word = 8'h0C;
		16'h74E: out_word = 8'h2A;
		16'h74F: out_word = 8'h4B;
		16'h750: out_word = 8'h5C;
		16'h751: out_word = 8'hED;
		16'h752: out_word = 8'h52;
		16'h753: out_word = 8'hDD;
		16'h754: out_word = 8'h75;
		16'h755: out_word = 8'h0F;
		16'h756: out_word = 8'hDD;
		16'h757: out_word = 8'h74;
		16'h758: out_word = 8'h10;
		16'h759: out_word = 8'hEB;
		16'h75A: out_word = 8'h3A;
		16'h75B: out_word = 8'h74;
		16'h75C: out_word = 8'h5C;
		16'h75D: out_word = 8'hA7;
		16'h75E: out_word = 8'hCA;
		16'h75F: out_word = 8'h70;
		16'h760: out_word = 8'h09;
		16'h761: out_word = 8'hE5;
		16'h762: out_word = 8'h01;
		16'h763: out_word = 8'h11;
		16'h764: out_word = 8'h00;
		16'h765: out_word = 8'hDD;
		16'h766: out_word = 8'h09;
		16'h767: out_word = 8'hDD;
		16'h768: out_word = 8'hE5;
		16'h769: out_word = 8'h11;
		16'h76A: out_word = 8'h11;
		16'h76B: out_word = 8'h00;
		16'h76C: out_word = 8'hAF;
		16'h76D: out_word = 8'h37;
		16'h76E: out_word = 8'hCD;
		16'h76F: out_word = 8'h56;
		16'h770: out_word = 8'h05;
		16'h771: out_word = 8'hDD;
		16'h772: out_word = 8'hE1;
		16'h773: out_word = 8'h30;
		16'h774: out_word = 8'hF2;
		16'h775: out_word = 8'h3E;
		16'h776: out_word = 8'hFE;
		16'h777: out_word = 8'hCD;
		16'h778: out_word = 8'h01;
		16'h779: out_word = 8'h16;
		16'h77A: out_word = 8'hFD;
		16'h77B: out_word = 8'h36;
		16'h77C: out_word = 8'h52;
		16'h77D: out_word = 8'h03;
		16'h77E: out_word = 8'h0E;
		16'h77F: out_word = 8'h80;
		16'h780: out_word = 8'hDD;
		16'h781: out_word = 8'h7E;
		16'h782: out_word = 8'h00;
		16'h783: out_word = 8'hDD;
		16'h784: out_word = 8'hBE;
		16'h785: out_word = 8'hEF;
		16'h786: out_word = 8'h20;
		16'h787: out_word = 8'h02;
		16'h788: out_word = 8'h0E;
		16'h789: out_word = 8'hF6;
		16'h78A: out_word = 8'hFE;
		16'h78B: out_word = 8'h04;
		16'h78C: out_word = 8'h30;
		16'h78D: out_word = 8'hD9;
		16'h78E: out_word = 8'h11;
		16'h78F: out_word = 8'hC0;
		16'h790: out_word = 8'h09;
		16'h791: out_word = 8'hC5;
		16'h792: out_word = 8'hCD;
		16'h793: out_word = 8'h0A;
		16'h794: out_word = 8'h0C;
		16'h795: out_word = 8'hC1;
		16'h796: out_word = 8'hDD;
		16'h797: out_word = 8'hE5;
		16'h798: out_word = 8'hD1;
		16'h799: out_word = 8'h21;
		16'h79A: out_word = 8'hF0;
		16'h79B: out_word = 8'hFF;
		16'h79C: out_word = 8'h19;
		16'h79D: out_word = 8'h06;
		16'h79E: out_word = 8'h0A;
		16'h79F: out_word = 8'h7E;
		16'h7A0: out_word = 8'h3C;
		16'h7A1: out_word = 8'h20;
		16'h7A2: out_word = 8'h03;
		16'h7A3: out_word = 8'h79;
		16'h7A4: out_word = 8'h80;
		16'h7A5: out_word = 8'h4F;
		16'h7A6: out_word = 8'h13;
		16'h7A7: out_word = 8'h1A;
		16'h7A8: out_word = 8'hBE;
		16'h7A9: out_word = 8'h23;
		16'h7AA: out_word = 8'h20;
		16'h7AB: out_word = 8'h01;
		16'h7AC: out_word = 8'h0C;
		16'h7AD: out_word = 8'hD7;
		16'h7AE: out_word = 8'h10;
		16'h7AF: out_word = 8'hF6;
		16'h7B0: out_word = 8'hCB;
		16'h7B1: out_word = 8'h79;
		16'h7B2: out_word = 8'h20;
		16'h7B3: out_word = 8'hB3;
		16'h7B4: out_word = 8'h3E;
		16'h7B5: out_word = 8'h0D;
		16'h7B6: out_word = 8'hD7;
		16'h7B7: out_word = 8'hE1;
		16'h7B8: out_word = 8'hDD;
		16'h7B9: out_word = 8'h7E;
		16'h7BA: out_word = 8'h00;
		16'h7BB: out_word = 8'hFE;
		16'h7BC: out_word = 8'h03;
		16'h7BD: out_word = 8'h28;
		16'h7BE: out_word = 8'h0C;
		16'h7BF: out_word = 8'h3A;
		16'h7C0: out_word = 8'h74;
		16'h7C1: out_word = 8'h5C;
		16'h7C2: out_word = 8'h3D;
		16'h7C3: out_word = 8'hCA;
		16'h7C4: out_word = 8'h08;
		16'h7C5: out_word = 8'h08;
		16'h7C6: out_word = 8'hFE;
		16'h7C7: out_word = 8'h02;
		16'h7C8: out_word = 8'hCA;
		16'h7C9: out_word = 8'hB6;
		16'h7CA: out_word = 8'h08;
		16'h7CB: out_word = 8'hE5;
		16'h7CC: out_word = 8'hDD;
		16'h7CD: out_word = 8'h6E;
		16'h7CE: out_word = 8'hFA;
		16'h7CF: out_word = 8'hDD;
		16'h7D0: out_word = 8'h66;
		16'h7D1: out_word = 8'hFB;
		16'h7D2: out_word = 8'hDD;
		16'h7D3: out_word = 8'h5E;
		16'h7D4: out_word = 8'h0B;
		16'h7D5: out_word = 8'hDD;
		16'h7D6: out_word = 8'h56;
		16'h7D7: out_word = 8'h0C;
		16'h7D8: out_word = 8'h7C;
		16'h7D9: out_word = 8'hB5;
		16'h7DA: out_word = 8'h28;
		16'h7DB: out_word = 8'h0D;
		16'h7DC: out_word = 8'hED;
		16'h7DD: out_word = 8'h52;
		16'h7DE: out_word = 8'h38;
		16'h7DF: out_word = 8'h26;
		16'h7E0: out_word = 8'h28;
		16'h7E1: out_word = 8'h07;
		16'h7E2: out_word = 8'hDD;
		16'h7E3: out_word = 8'h7E;
		16'h7E4: out_word = 8'h00;
		16'h7E5: out_word = 8'hFE;
		16'h7E6: out_word = 8'h03;
		16'h7E7: out_word = 8'h20;
		16'h7E8: out_word = 8'h1D;
		16'h7E9: out_word = 8'hE1;
		16'h7EA: out_word = 8'h7C;
		16'h7EB: out_word = 8'hB5;
		16'h7EC: out_word = 8'h20;
		16'h7ED: out_word = 8'h06;
		16'h7EE: out_word = 8'hDD;
		16'h7EF: out_word = 8'h6E;
		16'h7F0: out_word = 8'h0D;
		16'h7F1: out_word = 8'hDD;
		16'h7F2: out_word = 8'h66;
		16'h7F3: out_word = 8'h0E;
		16'h7F4: out_word = 8'hE5;
		16'h7F5: out_word = 8'hDD;
		16'h7F6: out_word = 8'hE1;
		16'h7F7: out_word = 8'h3A;
		16'h7F8: out_word = 8'h74;
		16'h7F9: out_word = 8'h5C;
		16'h7FA: out_word = 8'hFE;
		16'h7FB: out_word = 8'h02;
		16'h7FC: out_word = 8'h37;
		16'h7FD: out_word = 8'h20;
		16'h7FE: out_word = 8'h01;
		16'h7FF: out_word = 8'hA7;
		16'h800: out_word = 8'h3E;
		16'h801: out_word = 8'hFF;
		16'h802: out_word = 8'hCD;
		16'h803: out_word = 8'h56;
		16'h804: out_word = 8'h05;
		16'h805: out_word = 8'hD8;
		16'h806: out_word = 8'hCF;
		16'h807: out_word = 8'h1A;
		16'h808: out_word = 8'hDD;
		16'h809: out_word = 8'h5E;
		16'h80A: out_word = 8'h0B;
		16'h80B: out_word = 8'hDD;
		16'h80C: out_word = 8'h56;
		16'h80D: out_word = 8'h0C;
		16'h80E: out_word = 8'hE5;
		16'h80F: out_word = 8'h7C;
		16'h810: out_word = 8'hB5;
		16'h811: out_word = 8'h20;
		16'h812: out_word = 8'h06;
		16'h813: out_word = 8'h13;
		16'h814: out_word = 8'h13;
		16'h815: out_word = 8'h13;
		16'h816: out_word = 8'hEB;
		16'h817: out_word = 8'h18;
		16'h818: out_word = 8'h0C;
		16'h819: out_word = 8'hDD;
		16'h81A: out_word = 8'h6E;
		16'h81B: out_word = 8'hFA;
		16'h81C: out_word = 8'hDD;
		16'h81D: out_word = 8'h66;
		16'h81E: out_word = 8'hFB;
		16'h81F: out_word = 8'hEB;
		16'h820: out_word = 8'h37;
		16'h821: out_word = 8'hED;
		16'h822: out_word = 8'h52;
		16'h823: out_word = 8'h38;
		16'h824: out_word = 8'h09;
		16'h825: out_word = 8'h11;
		16'h826: out_word = 8'h05;
		16'h827: out_word = 8'h00;
		16'h828: out_word = 8'h19;
		16'h829: out_word = 8'h44;
		16'h82A: out_word = 8'h4D;
		16'h82B: out_word = 8'hCD;
		16'h82C: out_word = 8'h05;
		16'h82D: out_word = 8'h1F;
		16'h82E: out_word = 8'hE1;
		16'h82F: out_word = 8'hDD;
		16'h830: out_word = 8'h7E;
		16'h831: out_word = 8'h00;
		16'h832: out_word = 8'hA7;
		16'h833: out_word = 8'h28;
		16'h834: out_word = 8'h3E;
		16'h835: out_word = 8'h7C;
		16'h836: out_word = 8'hB5;
		16'h837: out_word = 8'h28;
		16'h838: out_word = 8'h13;
		16'h839: out_word = 8'h2B;
		16'h83A: out_word = 8'h46;
		16'h83B: out_word = 8'h2B;
		16'h83C: out_word = 8'h4E;
		16'h83D: out_word = 8'h2B;
		16'h83E: out_word = 8'h03;
		16'h83F: out_word = 8'h03;
		16'h840: out_word = 8'h03;
		16'h841: out_word = 8'hDD;
		16'h842: out_word = 8'h22;
		16'h843: out_word = 8'h5F;
		16'h844: out_word = 8'h5C;
		16'h845: out_word = 8'hCD;
		16'h846: out_word = 8'hE8;
		16'h847: out_word = 8'h19;
		16'h848: out_word = 8'hDD;
		16'h849: out_word = 8'h2A;
		16'h84A: out_word = 8'h5F;
		16'h84B: out_word = 8'h5C;
		16'h84C: out_word = 8'h2A;
		16'h84D: out_word = 8'h59;
		16'h84E: out_word = 8'h5C;
		16'h84F: out_word = 8'h2B;
		16'h850: out_word = 8'hDD;
		16'h851: out_word = 8'h4E;
		16'h852: out_word = 8'h0B;
		16'h853: out_word = 8'hDD;
		16'h854: out_word = 8'h46;
		16'h855: out_word = 8'h0C;
		16'h856: out_word = 8'hC5;
		16'h857: out_word = 8'h03;
		16'h858: out_word = 8'h03;
		16'h859: out_word = 8'h03;
		16'h85A: out_word = 8'hDD;
		16'h85B: out_word = 8'h7E;
		16'h85C: out_word = 8'hFD;
		16'h85D: out_word = 8'hF5;
		16'h85E: out_word = 8'hCD;
		16'h85F: out_word = 8'h55;
		16'h860: out_word = 8'h16;
		16'h861: out_word = 8'h23;
		16'h862: out_word = 8'hF1;
		16'h863: out_word = 8'h77;
		16'h864: out_word = 8'hD1;
		16'h865: out_word = 8'h23;
		16'h866: out_word = 8'h73;
		16'h867: out_word = 8'h23;
		16'h868: out_word = 8'h72;
		16'h869: out_word = 8'h23;
		16'h86A: out_word = 8'hE5;
		16'h86B: out_word = 8'hDD;
		16'h86C: out_word = 8'hE1;
		16'h86D: out_word = 8'h37;
		16'h86E: out_word = 8'h3E;
		16'h86F: out_word = 8'hFF;
		16'h870: out_word = 8'hC3;
		16'h871: out_word = 8'h02;
		16'h872: out_word = 8'h08;
		16'h873: out_word = 8'hEB;
		16'h874: out_word = 8'h2A;
		16'h875: out_word = 8'h59;
		16'h876: out_word = 8'h5C;
		16'h877: out_word = 8'h2B;
		16'h878: out_word = 8'hDD;
		16'h879: out_word = 8'h22;
		16'h87A: out_word = 8'h5F;
		16'h87B: out_word = 8'h5C;
		16'h87C: out_word = 8'hDD;
		16'h87D: out_word = 8'h4E;
		16'h87E: out_word = 8'h0B;
		16'h87F: out_word = 8'hDD;
		16'h880: out_word = 8'h46;
		16'h881: out_word = 8'h0C;
		16'h882: out_word = 8'hC5;
		16'h883: out_word = 8'hCD;
		16'h884: out_word = 8'hE5;
		16'h885: out_word = 8'h19;
		16'h886: out_word = 8'hC1;
		16'h887: out_word = 8'hE5;
		16'h888: out_word = 8'hC5;
		16'h889: out_word = 8'hCD;
		16'h88A: out_word = 8'h55;
		16'h88B: out_word = 8'h16;
		16'h88C: out_word = 8'hDD;
		16'h88D: out_word = 8'h2A;
		16'h88E: out_word = 8'h5F;
		16'h88F: out_word = 8'h5C;
		16'h890: out_word = 8'h23;
		16'h891: out_word = 8'hDD;
		16'h892: out_word = 8'h4E;
		16'h893: out_word = 8'h0F;
		16'h894: out_word = 8'hDD;
		16'h895: out_word = 8'h46;
		16'h896: out_word = 8'h10;
		16'h897: out_word = 8'h09;
		16'h898: out_word = 8'h22;
		16'h899: out_word = 8'h4B;
		16'h89A: out_word = 8'h5C;
		16'h89B: out_word = 8'hDD;
		16'h89C: out_word = 8'h66;
		16'h89D: out_word = 8'h0E;
		16'h89E: out_word = 8'h7C;
		16'h89F: out_word = 8'hE6;
		16'h8A0: out_word = 8'hC0;
		16'h8A1: out_word = 8'h20;
		16'h8A2: out_word = 8'h0A;
		16'h8A3: out_word = 8'hDD;
		16'h8A4: out_word = 8'h6E;
		16'h8A5: out_word = 8'h0D;
		16'h8A6: out_word = 8'h22;
		16'h8A7: out_word = 8'h42;
		16'h8A8: out_word = 8'h5C;
		16'h8A9: out_word = 8'hFD;
		16'h8AA: out_word = 8'h36;
		16'h8AB: out_word = 8'h0A;
		16'h8AC: out_word = 8'h00;
		16'h8AD: out_word = 8'hD1;
		16'h8AE: out_word = 8'hDD;
		16'h8AF: out_word = 8'hE1;
		16'h8B0: out_word = 8'h37;
		16'h8B1: out_word = 8'h3E;
		16'h8B2: out_word = 8'hFF;
		16'h8B3: out_word = 8'hC3;
		16'h8B4: out_word = 8'h02;
		16'h8B5: out_word = 8'h08;
		16'h8B6: out_word = 8'hDD;
		16'h8B7: out_word = 8'h4E;
		16'h8B8: out_word = 8'h0B;
		16'h8B9: out_word = 8'hDD;
		16'h8BA: out_word = 8'h46;
		16'h8BB: out_word = 8'h0C;
		16'h8BC: out_word = 8'hC5;
		16'h8BD: out_word = 8'h03;
		16'h8BE: out_word = 8'hF7;
		16'h8BF: out_word = 8'h36;
		16'h8C0: out_word = 8'h80;
		16'h8C1: out_word = 8'hEB;
		16'h8C2: out_word = 8'hD1;
		16'h8C3: out_word = 8'hE5;
		16'h8C4: out_word = 8'hE5;
		16'h8C5: out_word = 8'hDD;
		16'h8C6: out_word = 8'hE1;
		16'h8C7: out_word = 8'h37;
		16'h8C8: out_word = 8'h3E;
		16'h8C9: out_word = 8'hFF;
		16'h8CA: out_word = 8'hCD;
		16'h8CB: out_word = 8'h02;
		16'h8CC: out_word = 8'h08;
		16'h8CD: out_word = 8'hE1;
		16'h8CE: out_word = 8'hED;
		16'h8CF: out_word = 8'h5B;
		16'h8D0: out_word = 8'h53;
		16'h8D1: out_word = 8'h5C;
		16'h8D2: out_word = 8'h7E;
		16'h8D3: out_word = 8'hE6;
		16'h8D4: out_word = 8'hC0;
		16'h8D5: out_word = 8'h20;
		16'h8D6: out_word = 8'h19;
		16'h8D7: out_word = 8'h1A;
		16'h8D8: out_word = 8'h13;
		16'h8D9: out_word = 8'hBE;
		16'h8DA: out_word = 8'h23;
		16'h8DB: out_word = 8'h20;
		16'h8DC: out_word = 8'h02;
		16'h8DD: out_word = 8'h1A;
		16'h8DE: out_word = 8'hBE;
		16'h8DF: out_word = 8'h1B;
		16'h8E0: out_word = 8'h2B;
		16'h8E1: out_word = 8'h30;
		16'h8E2: out_word = 8'h08;
		16'h8E3: out_word = 8'hE5;
		16'h8E4: out_word = 8'hEB;
		16'h8E5: out_word = 8'hCD;
		16'h8E6: out_word = 8'hB8;
		16'h8E7: out_word = 8'h19;
		16'h8E8: out_word = 8'hE1;
		16'h8E9: out_word = 8'h18;
		16'h8EA: out_word = 8'hEC;
		16'h8EB: out_word = 8'hCD;
		16'h8EC: out_word = 8'h2C;
		16'h8ED: out_word = 8'h09;
		16'h8EE: out_word = 8'h18;
		16'h8EF: out_word = 8'hE2;
		16'h8F0: out_word = 8'h7E;
		16'h8F1: out_word = 8'h4F;
		16'h8F2: out_word = 8'hFE;
		16'h8F3: out_word = 8'h80;
		16'h8F4: out_word = 8'hC8;
		16'h8F5: out_word = 8'hE5;
		16'h8F6: out_word = 8'h2A;
		16'h8F7: out_word = 8'h4B;
		16'h8F8: out_word = 8'h5C;
		16'h8F9: out_word = 8'h7E;
		16'h8FA: out_word = 8'hFE;
		16'h8FB: out_word = 8'h80;
		16'h8FC: out_word = 8'h28;
		16'h8FD: out_word = 8'h25;
		16'h8FE: out_word = 8'hB9;
		16'h8FF: out_word = 8'h28;
		16'h900: out_word = 8'h08;
		16'h901: out_word = 8'hC5;
		16'h902: out_word = 8'hCD;
		16'h903: out_word = 8'hB8;
		16'h904: out_word = 8'h19;
		16'h905: out_word = 8'hC1;
		16'h906: out_word = 8'hEB;
		16'h907: out_word = 8'h18;
		16'h908: out_word = 8'hF0;
		16'h909: out_word = 8'hE6;
		16'h90A: out_word = 8'hE0;
		16'h90B: out_word = 8'hFE;
		16'h90C: out_word = 8'hA0;
		16'h90D: out_word = 8'h20;
		16'h90E: out_word = 8'h12;
		16'h90F: out_word = 8'hD1;
		16'h910: out_word = 8'hD5;
		16'h911: out_word = 8'hE5;
		16'h912: out_word = 8'h23;
		16'h913: out_word = 8'h13;
		16'h914: out_word = 8'h1A;
		16'h915: out_word = 8'hBE;
		16'h916: out_word = 8'h20;
		16'h917: out_word = 8'h06;
		16'h918: out_word = 8'h17;
		16'h919: out_word = 8'h30;
		16'h91A: out_word = 8'hF7;
		16'h91B: out_word = 8'hE1;
		16'h91C: out_word = 8'h18;
		16'h91D: out_word = 8'h03;
		16'h91E: out_word = 8'hE1;
		16'h91F: out_word = 8'h18;
		16'h920: out_word = 8'hE0;
		16'h921: out_word = 8'h3E;
		16'h922: out_word = 8'hFF;
		16'h923: out_word = 8'hD1;
		16'h924: out_word = 8'hEB;
		16'h925: out_word = 8'h3C;
		16'h926: out_word = 8'h37;
		16'h927: out_word = 8'hCD;
		16'h928: out_word = 8'h2C;
		16'h929: out_word = 8'h09;
		16'h92A: out_word = 8'h18;
		16'h92B: out_word = 8'hC4;
		16'h92C: out_word = 8'h20;
		16'h92D: out_word = 8'h10;
		16'h92E: out_word = 8'h08;
		16'h92F: out_word = 8'h22;
		16'h930: out_word = 8'h5F;
		16'h931: out_word = 8'h5C;
		16'h932: out_word = 8'hEB;
		16'h933: out_word = 8'hCD;
		16'h934: out_word = 8'hB8;
		16'h935: out_word = 8'h19;
		16'h936: out_word = 8'hCD;
		16'h937: out_word = 8'hE8;
		16'h938: out_word = 8'h19;
		16'h939: out_word = 8'hEB;
		16'h93A: out_word = 8'h2A;
		16'h93B: out_word = 8'h5F;
		16'h93C: out_word = 8'h5C;
		16'h93D: out_word = 8'h08;
		16'h93E: out_word = 8'h08;
		16'h93F: out_word = 8'hD5;
		16'h940: out_word = 8'hCD;
		16'h941: out_word = 8'hB8;
		16'h942: out_word = 8'h19;
		16'h943: out_word = 8'h22;
		16'h944: out_word = 8'h5F;
		16'h945: out_word = 8'h5C;
		16'h946: out_word = 8'h2A;
		16'h947: out_word = 8'h53;
		16'h948: out_word = 8'h5C;
		16'h949: out_word = 8'hE3;
		16'h94A: out_word = 8'hC5;
		16'h94B: out_word = 8'h08;
		16'h94C: out_word = 8'h38;
		16'h94D: out_word = 8'h07;
		16'h94E: out_word = 8'h2B;
		16'h94F: out_word = 8'hCD;
		16'h950: out_word = 8'h55;
		16'h951: out_word = 8'h16;
		16'h952: out_word = 8'h23;
		16'h953: out_word = 8'h18;
		16'h954: out_word = 8'h03;
		16'h955: out_word = 8'hCD;
		16'h956: out_word = 8'h55;
		16'h957: out_word = 8'h16;
		16'h958: out_word = 8'h23;
		16'h959: out_word = 8'hC1;
		16'h95A: out_word = 8'hD1;
		16'h95B: out_word = 8'hED;
		16'h95C: out_word = 8'h53;
		16'h95D: out_word = 8'h53;
		16'h95E: out_word = 8'h5C;
		16'h95F: out_word = 8'hED;
		16'h960: out_word = 8'h5B;
		16'h961: out_word = 8'h5F;
		16'h962: out_word = 8'h5C;
		16'h963: out_word = 8'hC5;
		16'h964: out_word = 8'hD5;
		16'h965: out_word = 8'hEB;
		16'h966: out_word = 8'hED;
		16'h967: out_word = 8'hB0;
		16'h968: out_word = 8'hE1;
		16'h969: out_word = 8'hC1;
		16'h96A: out_word = 8'hD5;
		16'h96B: out_word = 8'hCD;
		16'h96C: out_word = 8'hE8;
		16'h96D: out_word = 8'h19;
		16'h96E: out_word = 8'hD1;
		16'h96F: out_word = 8'hC9;
		16'h970: out_word = 8'hE5;
		16'h971: out_word = 8'h3E;
		16'h972: out_word = 8'hFD;
		16'h973: out_word = 8'hCD;
		16'h974: out_word = 8'h01;
		16'h975: out_word = 8'h16;
		16'h976: out_word = 8'hAF;
		16'h977: out_word = 8'h11;
		16'h978: out_word = 8'hA1;
		16'h979: out_word = 8'h09;
		16'h97A: out_word = 8'hCD;
		16'h97B: out_word = 8'h0A;
		16'h97C: out_word = 8'h0C;
		16'h97D: out_word = 8'hFD;
		16'h97E: out_word = 8'hCB;
		16'h97F: out_word = 8'h02;
		16'h980: out_word = 8'hEE;
		16'h981: out_word = 8'hCD;
		16'h982: out_word = 8'hD4;
		16'h983: out_word = 8'h15;
		16'h984: out_word = 8'hDD;
		16'h985: out_word = 8'hE5;
		16'h986: out_word = 8'h11;
		16'h987: out_word = 8'h11;
		16'h988: out_word = 8'h00;
		16'h989: out_word = 8'hAF;
		16'h98A: out_word = 8'hCD;
		16'h98B: out_word = 8'hC2;
		16'h98C: out_word = 8'h04;
		16'h98D: out_word = 8'hDD;
		16'h98E: out_word = 8'hE1;
		16'h98F: out_word = 8'h06;
		16'h990: out_word = 8'h32;
		16'h991: out_word = 8'h76;
		16'h992: out_word = 8'h10;
		16'h993: out_word = 8'hFD;
		16'h994: out_word = 8'hDD;
		16'h995: out_word = 8'h5E;
		16'h996: out_word = 8'h0B;
		16'h997: out_word = 8'hDD;
		16'h998: out_word = 8'h56;
		16'h999: out_word = 8'h0C;
		16'h99A: out_word = 8'h3E;
		16'h99B: out_word = 8'hFF;
		16'h99C: out_word = 8'hDD;
		16'h99D: out_word = 8'hE1;
		16'h99E: out_word = 8'hC3;
		16'h99F: out_word = 8'hC2;
		16'h9A0: out_word = 8'h04;
		16'h9A1: out_word = 8'h80;
		16'h9A2: out_word = 8'h53;
		16'h9A3: out_word = 8'h74;
		16'h9A4: out_word = 8'h61;
		16'h9A5: out_word = 8'h72;
		16'h9A6: out_word = 8'h74;
		16'h9A7: out_word = 8'h20;
		16'h9A8: out_word = 8'h74;
		16'h9A9: out_word = 8'h61;
		16'h9AA: out_word = 8'h70;
		16'h9AB: out_word = 8'h65;
		16'h9AC: out_word = 8'h2C;
		16'h9AD: out_word = 8'h20;
		16'h9AE: out_word = 8'h74;
		16'h9AF: out_word = 8'h68;
		16'h9B0: out_word = 8'h65;
		16'h9B1: out_word = 8'h6E;
		16'h9B2: out_word = 8'h20;
		16'h9B3: out_word = 8'h70;
		16'h9B4: out_word = 8'h72;
		16'h9B5: out_word = 8'h65;
		16'h9B6: out_word = 8'h73;
		16'h9B7: out_word = 8'h73;
		16'h9B8: out_word = 8'h20;
		16'h9B9: out_word = 8'h61;
		16'h9BA: out_word = 8'h6E;
		16'h9BB: out_word = 8'h79;
		16'h9BC: out_word = 8'h20;
		16'h9BD: out_word = 8'h6B;
		16'h9BE: out_word = 8'h65;
		16'h9BF: out_word = 8'h79;
		16'h9C0: out_word = 8'hAE;
		16'h9C1: out_word = 8'h0D;
		16'h9C2: out_word = 8'h50;
		16'h9C3: out_word = 8'h72;
		16'h9C4: out_word = 8'h6F;
		16'h9C5: out_word = 8'h67;
		16'h9C6: out_word = 8'h72;
		16'h9C7: out_word = 8'h61;
		16'h9C8: out_word = 8'h6D;
		16'h9C9: out_word = 8'h3A;
		16'h9CA: out_word = 8'hA0;
		16'h9CB: out_word = 8'h0D;
		16'h9CC: out_word = 8'h4E;
		16'h9CD: out_word = 8'h75;
		16'h9CE: out_word = 8'h6D;
		16'h9CF: out_word = 8'h62;
		16'h9D0: out_word = 8'h65;
		16'h9D1: out_word = 8'h72;
		16'h9D2: out_word = 8'h20;
		16'h9D3: out_word = 8'h61;
		16'h9D4: out_word = 8'h72;
		16'h9D5: out_word = 8'h72;
		16'h9D6: out_word = 8'h61;
		16'h9D7: out_word = 8'h79;
		16'h9D8: out_word = 8'h3A;
		16'h9D9: out_word = 8'hA0;
		16'h9DA: out_word = 8'h0D;
		16'h9DB: out_word = 8'h43;
		16'h9DC: out_word = 8'h68;
		16'h9DD: out_word = 8'h61;
		16'h9DE: out_word = 8'h72;
		16'h9DF: out_word = 8'h61;
		16'h9E0: out_word = 8'h63;
		16'h9E1: out_word = 8'h74;
		16'h9E2: out_word = 8'h65;
		16'h9E3: out_word = 8'h72;
		16'h9E4: out_word = 8'h20;
		16'h9E5: out_word = 8'h61;
		16'h9E6: out_word = 8'h72;
		16'h9E7: out_word = 8'h72;
		16'h9E8: out_word = 8'h61;
		16'h9E9: out_word = 8'h79;
		16'h9EA: out_word = 8'h3A;
		16'h9EB: out_word = 8'hA0;
		16'h9EC: out_word = 8'h0D;
		16'h9ED: out_word = 8'h42;
		16'h9EE: out_word = 8'h79;
		16'h9EF: out_word = 8'h74;
		16'h9F0: out_word = 8'h65;
		16'h9F1: out_word = 8'h73;
		16'h9F2: out_word = 8'h3A;
		16'h9F3: out_word = 8'hA0;
		16'h9F4: out_word = 8'hCD;
		16'h9F5: out_word = 8'h03;
		16'h9F6: out_word = 8'h0B;
		16'h9F7: out_word = 8'hFE;
		16'h9F8: out_word = 8'h20;
		16'h9F9: out_word = 8'hD2;
		16'h9FA: out_word = 8'hD9;
		16'h9FB: out_word = 8'h0A;
		16'h9FC: out_word = 8'hFE;
		16'h9FD: out_word = 8'h06;
		16'h9FE: out_word = 8'h38;
		16'h9FF: out_word = 8'h69;
		16'hA00: out_word = 8'hFE;
		16'hA01: out_word = 8'h18;
		16'hA02: out_word = 8'h30;
		16'hA03: out_word = 8'h65;
		16'hA04: out_word = 8'h21;
		16'hA05: out_word = 8'h0B;
		16'hA06: out_word = 8'h0A;
		16'hA07: out_word = 8'h5F;
		16'hA08: out_word = 8'h16;
		16'hA09: out_word = 8'h00;
		16'hA0A: out_word = 8'h19;
		16'hA0B: out_word = 8'h5E;
		16'hA0C: out_word = 8'h19;
		16'hA0D: out_word = 8'hE5;
		16'hA0E: out_word = 8'hC3;
		16'hA0F: out_word = 8'h03;
		16'hA10: out_word = 8'h0B;
		16'hA11: out_word = 8'h4E;
		16'hA12: out_word = 8'h57;
		16'hA13: out_word = 8'h10;
		16'hA14: out_word = 8'h29;
		16'hA15: out_word = 8'h54;
		16'hA16: out_word = 8'h53;
		16'hA17: out_word = 8'h52;
		16'hA18: out_word = 8'h37;
		16'hA19: out_word = 8'h50;
		16'hA1A: out_word = 8'h4F;
		16'hA1B: out_word = 8'h5F;
		16'hA1C: out_word = 8'h5E;
		16'hA1D: out_word = 8'h5D;
		16'hA1E: out_word = 8'h5C;
		16'hA1F: out_word = 8'h5B;
		16'hA20: out_word = 8'h5A;
		16'hA21: out_word = 8'h54;
		16'hA22: out_word = 8'h53;
		16'hA23: out_word = 8'h0C;
		16'hA24: out_word = 8'h3E;
		16'hA25: out_word = 8'h22;
		16'hA26: out_word = 8'hB9;
		16'hA27: out_word = 8'h20;
		16'hA28: out_word = 8'h11;
		16'hA29: out_word = 8'hFD;
		16'hA2A: out_word = 8'hCB;
		16'hA2B: out_word = 8'h01;
		16'hA2C: out_word = 8'h4E;
		16'hA2D: out_word = 8'h20;
		16'hA2E: out_word = 8'h09;
		16'hA2F: out_word = 8'h04;
		16'hA30: out_word = 8'h0E;
		16'hA31: out_word = 8'h02;
		16'hA32: out_word = 8'h3E;
		16'hA33: out_word = 8'h18;
		16'hA34: out_word = 8'hB8;
		16'hA35: out_word = 8'h20;
		16'hA36: out_word = 8'h03;
		16'hA37: out_word = 8'h05;
		16'hA38: out_word = 8'h0E;
		16'hA39: out_word = 8'h21;
		16'hA3A: out_word = 8'hC3;
		16'hA3B: out_word = 8'hD9;
		16'hA3C: out_word = 8'h0D;
		16'hA3D: out_word = 8'h3A;
		16'hA3E: out_word = 8'h91;
		16'hA3F: out_word = 8'h5C;
		16'hA40: out_word = 8'hF5;
		16'hA41: out_word = 8'hFD;
		16'hA42: out_word = 8'h36;
		16'hA43: out_word = 8'h57;
		16'hA44: out_word = 8'h01;
		16'hA45: out_word = 8'h3E;
		16'hA46: out_word = 8'h20;
		16'hA47: out_word = 8'hCD;
		16'hA48: out_word = 8'h65;
		16'hA49: out_word = 8'h0B;
		16'hA4A: out_word = 8'hF1;
		16'hA4B: out_word = 8'h32;
		16'hA4C: out_word = 8'h91;
		16'hA4D: out_word = 8'h5C;
		16'hA4E: out_word = 8'hC9;
		16'hA4F: out_word = 8'hFD;
		16'hA50: out_word = 8'hCB;
		16'hA51: out_word = 8'h01;
		16'hA52: out_word = 8'h4E;
		16'hA53: out_word = 8'hC2;
		16'hA54: out_word = 8'hCD;
		16'hA55: out_word = 8'h0E;
		16'hA56: out_word = 8'h0E;
		16'hA57: out_word = 8'h21;
		16'hA58: out_word = 8'hCD;
		16'hA59: out_word = 8'h55;
		16'hA5A: out_word = 8'h0C;
		16'hA5B: out_word = 8'h05;
		16'hA5C: out_word = 8'hC3;
		16'hA5D: out_word = 8'hD9;
		16'hA5E: out_word = 8'h0D;
		16'hA5F: out_word = 8'hCD;
		16'hA60: out_word = 8'h03;
		16'hA61: out_word = 8'h0B;
		16'hA62: out_word = 8'h79;
		16'hA63: out_word = 8'h3D;
		16'hA64: out_word = 8'h3D;
		16'hA65: out_word = 8'hE6;
		16'hA66: out_word = 8'h10;
		16'hA67: out_word = 8'h18;
		16'hA68: out_word = 8'h5A;
		16'hA69: out_word = 8'h3E;
		16'hA6A: out_word = 8'h3F;
		16'hA6B: out_word = 8'h18;
		16'hA6C: out_word = 8'h6C;
		16'hA6D: out_word = 8'h11;
		16'hA6E: out_word = 8'h87;
		16'hA6F: out_word = 8'h0A;
		16'hA70: out_word = 8'h32;
		16'hA71: out_word = 8'h0F;
		16'hA72: out_word = 8'h5C;
		16'hA73: out_word = 8'h18;
		16'hA74: out_word = 8'h0B;
		16'hA75: out_word = 8'h11;
		16'hA76: out_word = 8'h6D;
		16'hA77: out_word = 8'h0A;
		16'hA78: out_word = 8'h18;
		16'hA79: out_word = 8'h03;
		16'hA7A: out_word = 8'h11;
		16'hA7B: out_word = 8'h87;
		16'hA7C: out_word = 8'h0A;
		16'hA7D: out_word = 8'h32;
		16'hA7E: out_word = 8'h0E;
		16'hA7F: out_word = 8'h5C;
		16'hA80: out_word = 8'h2A;
		16'hA81: out_word = 8'h51;
		16'hA82: out_word = 8'h5C;
		16'hA83: out_word = 8'h73;
		16'hA84: out_word = 8'h23;
		16'hA85: out_word = 8'h72;
		16'hA86: out_word = 8'hC9;
		16'hA87: out_word = 8'h11;
		16'hA88: out_word = 8'hF4;
		16'hA89: out_word = 8'h09;
		16'hA8A: out_word = 8'hCD;
		16'hA8B: out_word = 8'h80;
		16'hA8C: out_word = 8'h0A;
		16'hA8D: out_word = 8'h2A;
		16'hA8E: out_word = 8'h0E;
		16'hA8F: out_word = 8'h5C;
		16'hA90: out_word = 8'h57;
		16'hA91: out_word = 8'h7D;
		16'hA92: out_word = 8'hFE;
		16'hA93: out_word = 8'h16;
		16'hA94: out_word = 8'hDA;
		16'hA95: out_word = 8'h11;
		16'hA96: out_word = 8'h22;
		16'hA97: out_word = 8'h20;
		16'hA98: out_word = 8'h29;
		16'hA99: out_word = 8'h44;
		16'hA9A: out_word = 8'h4A;
		16'hA9B: out_word = 8'h3E;
		16'hA9C: out_word = 8'h1F;
		16'hA9D: out_word = 8'h91;
		16'hA9E: out_word = 8'h38;
		16'hA9F: out_word = 8'h0C;
		16'hAA0: out_word = 8'hC6;
		16'hAA1: out_word = 8'h02;
		16'hAA2: out_word = 8'h4F;
		16'hAA3: out_word = 8'hFD;
		16'hAA4: out_word = 8'hCB;
		16'hAA5: out_word = 8'h01;
		16'hAA6: out_word = 8'h4E;
		16'hAA7: out_word = 8'h20;
		16'hAA8: out_word = 8'h16;
		16'hAA9: out_word = 8'h3E;
		16'hAAA: out_word = 8'h16;
		16'hAAB: out_word = 8'h90;
		16'hAAC: out_word = 8'hDA;
		16'hAAD: out_word = 8'h9F;
		16'hAAE: out_word = 8'h1E;
		16'hAAF: out_word = 8'h3C;
		16'hAB0: out_word = 8'h47;
		16'hAB1: out_word = 8'h04;
		16'hAB2: out_word = 8'hFD;
		16'hAB3: out_word = 8'hCB;
		16'hAB4: out_word = 8'h02;
		16'hAB5: out_word = 8'h46;
		16'hAB6: out_word = 8'hC2;
		16'hAB7: out_word = 8'h55;
		16'hAB8: out_word = 8'h0C;
		16'hAB9: out_word = 8'hFD;
		16'hABA: out_word = 8'hBE;
		16'hABB: out_word = 8'h31;
		16'hABC: out_word = 8'hDA;
		16'hABD: out_word = 8'h86;
		16'hABE: out_word = 8'h0C;
		16'hABF: out_word = 8'hC3;
		16'hAC0: out_word = 8'hD9;
		16'hAC1: out_word = 8'h0D;
		16'hAC2: out_word = 8'h7C;
		16'hAC3: out_word = 8'hCD;
		16'hAC4: out_word = 8'h03;
		16'hAC5: out_word = 8'h0B;
		16'hAC6: out_word = 8'h81;
		16'hAC7: out_word = 8'h3D;
		16'hAC8: out_word = 8'hE6;
		16'hAC9: out_word = 8'h1F;
		16'hACA: out_word = 8'hC8;
		16'hACB: out_word = 8'h57;
		16'hACC: out_word = 8'hFD;
		16'hACD: out_word = 8'hCB;
		16'hACE: out_word = 8'h01;
		16'hACF: out_word = 8'hC6;
		16'hAD0: out_word = 8'h3E;
		16'hAD1: out_word = 8'h20;
		16'hAD2: out_word = 8'hCD;
		16'hAD3: out_word = 8'h3B;
		16'hAD4: out_word = 8'h0C;
		16'hAD5: out_word = 8'h15;
		16'hAD6: out_word = 8'h20;
		16'hAD7: out_word = 8'hF8;
		16'hAD8: out_word = 8'hC9;
		16'hAD9: out_word = 8'hCD;
		16'hADA: out_word = 8'h24;
		16'hADB: out_word = 8'h0B;
		16'hADC: out_word = 8'hFD;
		16'hADD: out_word = 8'hCB;
		16'hADE: out_word = 8'h01;
		16'hADF: out_word = 8'h4E;
		16'hAE0: out_word = 8'h20;
		16'hAE1: out_word = 8'h1A;
		16'hAE2: out_word = 8'hFD;
		16'hAE3: out_word = 8'hCB;
		16'hAE4: out_word = 8'h02;
		16'hAE5: out_word = 8'h46;
		16'hAE6: out_word = 8'h20;
		16'hAE7: out_word = 8'h08;
		16'hAE8: out_word = 8'hED;
		16'hAE9: out_word = 8'h43;
		16'hAEA: out_word = 8'h88;
		16'hAEB: out_word = 8'h5C;
		16'hAEC: out_word = 8'h22;
		16'hAED: out_word = 8'h84;
		16'hAEE: out_word = 8'h5C;
		16'hAEF: out_word = 8'hC9;
		16'hAF0: out_word = 8'hED;
		16'hAF1: out_word = 8'h43;
		16'hAF2: out_word = 8'h8A;
		16'hAF3: out_word = 8'h5C;
		16'hAF4: out_word = 8'hED;
		16'hAF5: out_word = 8'h43;
		16'hAF6: out_word = 8'h82;
		16'hAF7: out_word = 8'h5C;
		16'hAF8: out_word = 8'h22;
		16'hAF9: out_word = 8'h86;
		16'hAFA: out_word = 8'h5C;
		16'hAFB: out_word = 8'hC9;
		16'hAFC: out_word = 8'hFD;
		16'hAFD: out_word = 8'h71;
		16'hAFE: out_word = 8'h45;
		16'hAFF: out_word = 8'h22;
		16'hB00: out_word = 8'h80;
		16'hB01: out_word = 8'h5C;
		16'hB02: out_word = 8'hC9;
		16'hB03: out_word = 8'hFD;
		16'hB04: out_word = 8'hCB;
		16'hB05: out_word = 8'h01;
		16'hB06: out_word = 8'h4E;
		16'hB07: out_word = 8'h20;
		16'hB08: out_word = 8'h14;
		16'hB09: out_word = 8'hED;
		16'hB0A: out_word = 8'h4B;
		16'hB0B: out_word = 8'h88;
		16'hB0C: out_word = 8'h5C;
		16'hB0D: out_word = 8'h2A;
		16'hB0E: out_word = 8'h84;
		16'hB0F: out_word = 8'h5C;
		16'hB10: out_word = 8'hFD;
		16'hB11: out_word = 8'hCB;
		16'hB12: out_word = 8'h02;
		16'hB13: out_word = 8'h46;
		16'hB14: out_word = 8'hC8;
		16'hB15: out_word = 8'hED;
		16'hB16: out_word = 8'h4B;
		16'hB17: out_word = 8'h8A;
		16'hB18: out_word = 8'h5C;
		16'hB19: out_word = 8'h2A;
		16'hB1A: out_word = 8'h86;
		16'hB1B: out_word = 8'h5C;
		16'hB1C: out_word = 8'hC9;
		16'hB1D: out_word = 8'hFD;
		16'hB1E: out_word = 8'h4E;
		16'hB1F: out_word = 8'h45;
		16'hB20: out_word = 8'h2A;
		16'hB21: out_word = 8'h80;
		16'hB22: out_word = 8'h5C;
		16'hB23: out_word = 8'hC9;
		16'hB24: out_word = 8'hFE;
		16'hB25: out_word = 8'h80;
		16'hB26: out_word = 8'h38;
		16'hB27: out_word = 8'h3D;
		16'hB28: out_word = 8'hFE;
		16'hB29: out_word = 8'h90;
		16'hB2A: out_word = 8'h30;
		16'hB2B: out_word = 8'h26;
		16'hB2C: out_word = 8'h47;
		16'hB2D: out_word = 8'hCD;
		16'hB2E: out_word = 8'h38;
		16'hB2F: out_word = 8'h0B;
		16'hB30: out_word = 8'hCD;
		16'hB31: out_word = 8'h03;
		16'hB32: out_word = 8'h0B;
		16'hB33: out_word = 8'h11;
		16'hB34: out_word = 8'h92;
		16'hB35: out_word = 8'h5C;
		16'hB36: out_word = 8'h18;
		16'hB37: out_word = 8'h47;
		16'hB38: out_word = 8'h21;
		16'hB39: out_word = 8'h92;
		16'hB3A: out_word = 8'h5C;
		16'hB3B: out_word = 8'hCD;
		16'hB3C: out_word = 8'h3E;
		16'hB3D: out_word = 8'h0B;
		16'hB3E: out_word = 8'hCB;
		16'hB3F: out_word = 8'h18;
		16'hB40: out_word = 8'h9F;
		16'hB41: out_word = 8'hE6;
		16'hB42: out_word = 8'h0F;
		16'hB43: out_word = 8'h4F;
		16'hB44: out_word = 8'hCB;
		16'hB45: out_word = 8'h18;
		16'hB46: out_word = 8'h9F;
		16'hB47: out_word = 8'hE6;
		16'hB48: out_word = 8'hF0;
		16'hB49: out_word = 8'hB1;
		16'hB4A: out_word = 8'h0E;
		16'hB4B: out_word = 8'h04;
		16'hB4C: out_word = 8'h77;
		16'hB4D: out_word = 8'h23;
		16'hB4E: out_word = 8'h0D;
		16'hB4F: out_word = 8'h20;
		16'hB50: out_word = 8'hFB;
		16'hB51: out_word = 8'hC9;
		16'hB52: out_word = 8'hC3;
		16'hB53: out_word = 8'h9F;
		16'hB54: out_word = 8'h3B;
		16'hB55: out_word = 8'h00;
		16'hB56: out_word = 8'hC6;
		16'hB57: out_word = 8'h15;
		16'hB58: out_word = 8'hC5;
		16'hB59: out_word = 8'hED;
		16'hB5A: out_word = 8'h4B;
		16'hB5B: out_word = 8'h7B;
		16'hB5C: out_word = 8'h5C;
		16'hB5D: out_word = 8'h18;
		16'hB5E: out_word = 8'h0B;
		16'hB5F: out_word = 8'hCD;
		16'hB60: out_word = 8'h10;
		16'hB61: out_word = 8'h0C;
		16'hB62: out_word = 8'hC3;
		16'hB63: out_word = 8'h03;
		16'hB64: out_word = 8'h0B;
		16'hB65: out_word = 8'hC5;
		16'hB66: out_word = 8'hED;
		16'hB67: out_word = 8'h4B;
		16'hB68: out_word = 8'h36;
		16'hB69: out_word = 8'h5C;
		16'hB6A: out_word = 8'hEB;
		16'hB6B: out_word = 8'h21;
		16'hB6C: out_word = 8'h3B;
		16'hB6D: out_word = 8'h5C;
		16'hB6E: out_word = 8'hCB;
		16'hB6F: out_word = 8'h86;
		16'hB70: out_word = 8'hFE;
		16'hB71: out_word = 8'h20;
		16'hB72: out_word = 8'h20;
		16'hB73: out_word = 8'h02;
		16'hB74: out_word = 8'hCB;
		16'hB75: out_word = 8'hC6;
		16'hB76: out_word = 8'h26;
		16'hB77: out_word = 8'h00;
		16'hB78: out_word = 8'h6F;
		16'hB79: out_word = 8'h29;
		16'hB7A: out_word = 8'h29;
		16'hB7B: out_word = 8'h29;
		16'hB7C: out_word = 8'h09;
		16'hB7D: out_word = 8'hC1;
		16'hB7E: out_word = 8'hEB;
		16'hB7F: out_word = 8'h79;
		16'hB80: out_word = 8'h3D;
		16'hB81: out_word = 8'h3E;
		16'hB82: out_word = 8'h21;
		16'hB83: out_word = 8'h20;
		16'hB84: out_word = 8'h0E;
		16'hB85: out_word = 8'h05;
		16'hB86: out_word = 8'h4F;
		16'hB87: out_word = 8'hFD;
		16'hB88: out_word = 8'hCB;
		16'hB89: out_word = 8'h01;
		16'hB8A: out_word = 8'h4E;
		16'hB8B: out_word = 8'h28;
		16'hB8C: out_word = 8'h06;
		16'hB8D: out_word = 8'hD5;
		16'hB8E: out_word = 8'hCD;
		16'hB8F: out_word = 8'hCD;
		16'hB90: out_word = 8'h0E;
		16'hB91: out_word = 8'hD1;
		16'hB92: out_word = 8'h79;
		16'hB93: out_word = 8'hB9;
		16'hB94: out_word = 8'hD5;
		16'hB95: out_word = 8'hCC;
		16'hB96: out_word = 8'h55;
		16'hB97: out_word = 8'h0C;
		16'hB98: out_word = 8'hD1;
		16'hB99: out_word = 8'hC5;
		16'hB9A: out_word = 8'hE5;
		16'hB9B: out_word = 8'h3A;
		16'hB9C: out_word = 8'h91;
		16'hB9D: out_word = 8'h5C;
		16'hB9E: out_word = 8'h06;
		16'hB9F: out_word = 8'hFF;
		16'hBA0: out_word = 8'h1F;
		16'hBA1: out_word = 8'h38;
		16'hBA2: out_word = 8'h01;
		16'hBA3: out_word = 8'h04;
		16'hBA4: out_word = 8'h1F;
		16'hBA5: out_word = 8'h1F;
		16'hBA6: out_word = 8'h9F;
		16'hBA7: out_word = 8'h4F;
		16'hBA8: out_word = 8'h3E;
		16'hBA9: out_word = 8'h08;
		16'hBAA: out_word = 8'hA7;
		16'hBAB: out_word = 8'hFD;
		16'hBAC: out_word = 8'hCB;
		16'hBAD: out_word = 8'h01;
		16'hBAE: out_word = 8'h4E;
		16'hBAF: out_word = 8'h28;
		16'hBB0: out_word = 8'h05;
		16'hBB1: out_word = 8'hFD;
		16'hBB2: out_word = 8'hCB;
		16'hBB3: out_word = 8'h30;
		16'hBB4: out_word = 8'hCE;
		16'hBB5: out_word = 8'h37;
		16'hBB6: out_word = 8'hEB;
		16'hBB7: out_word = 8'h08;
		16'hBB8: out_word = 8'h1A;
		16'hBB9: out_word = 8'hA0;
		16'hBBA: out_word = 8'hAE;
		16'hBBB: out_word = 8'hA9;
		16'hBBC: out_word = 8'h12;
		16'hBBD: out_word = 8'h08;
		16'hBBE: out_word = 8'h38;
		16'hBBF: out_word = 8'h13;
		16'hBC0: out_word = 8'h14;
		16'hBC1: out_word = 8'h23;
		16'hBC2: out_word = 8'h3D;
		16'hBC3: out_word = 8'h20;
		16'hBC4: out_word = 8'hF2;
		16'hBC5: out_word = 8'hEB;
		16'hBC6: out_word = 8'h25;
		16'hBC7: out_word = 8'hFD;
		16'hBC8: out_word = 8'hCB;
		16'hBC9: out_word = 8'h01;
		16'hBCA: out_word = 8'h4E;
		16'hBCB: out_word = 8'hCC;
		16'hBCC: out_word = 8'hDB;
		16'hBCD: out_word = 8'h0B;
		16'hBCE: out_word = 8'hE1;
		16'hBCF: out_word = 8'hC1;
		16'hBD0: out_word = 8'h0D;
		16'hBD1: out_word = 8'h23;
		16'hBD2: out_word = 8'hC9;
		16'hBD3: out_word = 8'h08;
		16'hBD4: out_word = 8'h3E;
		16'hBD5: out_word = 8'h20;
		16'hBD6: out_word = 8'h83;
		16'hBD7: out_word = 8'h5F;
		16'hBD8: out_word = 8'h08;
		16'hBD9: out_word = 8'h18;
		16'hBDA: out_word = 8'hE6;
		16'hBDB: out_word = 8'h7C;
		16'hBDC: out_word = 8'h0F;
		16'hBDD: out_word = 8'h0F;
		16'hBDE: out_word = 8'h0F;
		16'hBDF: out_word = 8'hE6;
		16'hBE0: out_word = 8'h03;
		16'hBE1: out_word = 8'hF6;
		16'hBE2: out_word = 8'h58;
		16'hBE3: out_word = 8'h67;
		16'hBE4: out_word = 8'hED;
		16'hBE5: out_word = 8'h5B;
		16'hBE6: out_word = 8'h8F;
		16'hBE7: out_word = 8'h5C;
		16'hBE8: out_word = 8'h7E;
		16'hBE9: out_word = 8'hAB;
		16'hBEA: out_word = 8'hA2;
		16'hBEB: out_word = 8'hAB;
		16'hBEC: out_word = 8'hFD;
		16'hBED: out_word = 8'hCB;
		16'hBEE: out_word = 8'h57;
		16'hBEF: out_word = 8'h76;
		16'hBF0: out_word = 8'h28;
		16'hBF1: out_word = 8'h08;
		16'hBF2: out_word = 8'hE6;
		16'hBF3: out_word = 8'hC7;
		16'hBF4: out_word = 8'hCB;
		16'hBF5: out_word = 8'h57;
		16'hBF6: out_word = 8'h20;
		16'hBF7: out_word = 8'h02;
		16'hBF8: out_word = 8'hEE;
		16'hBF9: out_word = 8'h38;
		16'hBFA: out_word = 8'hFD;
		16'hBFB: out_word = 8'hCB;
		16'hBFC: out_word = 8'h57;
		16'hBFD: out_word = 8'h66;
		16'hBFE: out_word = 8'h28;
		16'hBFF: out_word = 8'h08;
		16'hC00: out_word = 8'hE6;
		16'hC01: out_word = 8'hF8;
		16'hC02: out_word = 8'hCB;
		16'hC03: out_word = 8'h6F;
		16'hC04: out_word = 8'h20;
		16'hC05: out_word = 8'h02;
		16'hC06: out_word = 8'hEE;
		16'hC07: out_word = 8'h07;
		16'hC08: out_word = 8'h77;
		16'hC09: out_word = 8'hC9;
		16'hC0A: out_word = 8'hE5;
		16'hC0B: out_word = 8'h26;
		16'hC0C: out_word = 8'h00;
		16'hC0D: out_word = 8'hE3;
		16'hC0E: out_word = 8'h18;
		16'hC0F: out_word = 8'h04;
		16'hC10: out_word = 8'h11;
		16'hC11: out_word = 8'h95;
		16'hC12: out_word = 8'h00;
		16'hC13: out_word = 8'hF5;
		16'hC14: out_word = 8'hCD;
		16'hC15: out_word = 8'h41;
		16'hC16: out_word = 8'h0C;
		16'hC17: out_word = 8'h38;
		16'hC18: out_word = 8'h09;
		16'hC19: out_word = 8'h3E;
		16'hC1A: out_word = 8'h20;
		16'hC1B: out_word = 8'hFD;
		16'hC1C: out_word = 8'hCB;
		16'hC1D: out_word = 8'h01;
		16'hC1E: out_word = 8'h46;
		16'hC1F: out_word = 8'hCC;
		16'hC20: out_word = 8'h3B;
		16'hC21: out_word = 8'h0C;
		16'hC22: out_word = 8'h1A;
		16'hC23: out_word = 8'hE6;
		16'hC24: out_word = 8'h7F;
		16'hC25: out_word = 8'hCD;
		16'hC26: out_word = 8'h3B;
		16'hC27: out_word = 8'h0C;
		16'hC28: out_word = 8'h1A;
		16'hC29: out_word = 8'h13;
		16'hC2A: out_word = 8'h87;
		16'hC2B: out_word = 8'h30;
		16'hC2C: out_word = 8'hF5;
		16'hC2D: out_word = 8'hD1;
		16'hC2E: out_word = 8'hFE;
		16'hC2F: out_word = 8'h48;
		16'hC30: out_word = 8'h28;
		16'hC31: out_word = 8'h03;
		16'hC32: out_word = 8'hFE;
		16'hC33: out_word = 8'h82;
		16'hC34: out_word = 8'hD8;
		16'hC35: out_word = 8'h7A;
		16'hC36: out_word = 8'hFE;
		16'hC37: out_word = 8'h03;
		16'hC38: out_word = 8'hD8;
		16'hC39: out_word = 8'h3E;
		16'hC3A: out_word = 8'h20;
		16'hC3B: out_word = 8'hD5;
		16'hC3C: out_word = 8'hD9;
		16'hC3D: out_word = 8'hD7;
		16'hC3E: out_word = 8'hD9;
		16'hC3F: out_word = 8'hD1;
		16'hC40: out_word = 8'hC9;
		16'hC41: out_word = 8'hF5;
		16'hC42: out_word = 8'hEB;
		16'hC43: out_word = 8'h3C;
		16'hC44: out_word = 8'hCB;
		16'hC45: out_word = 8'h7E;
		16'hC46: out_word = 8'h23;
		16'hC47: out_word = 8'h28;
		16'hC48: out_word = 8'hFB;
		16'hC49: out_word = 8'h3D;
		16'hC4A: out_word = 8'h20;
		16'hC4B: out_word = 8'hF8;
		16'hC4C: out_word = 8'hEB;
		16'hC4D: out_word = 8'hF1;
		16'hC4E: out_word = 8'hFE;
		16'hC4F: out_word = 8'h20;
		16'hC50: out_word = 8'hD8;
		16'hC51: out_word = 8'h1A;
		16'hC52: out_word = 8'hD6;
		16'hC53: out_word = 8'h41;
		16'hC54: out_word = 8'hC9;
		16'hC55: out_word = 8'hFD;
		16'hC56: out_word = 8'hCB;
		16'hC57: out_word = 8'h01;
		16'hC58: out_word = 8'h4E;
		16'hC59: out_word = 8'hC0;
		16'hC5A: out_word = 8'h11;
		16'hC5B: out_word = 8'hD9;
		16'hC5C: out_word = 8'h0D;
		16'hC5D: out_word = 8'hD5;
		16'hC5E: out_word = 8'h78;
		16'hC5F: out_word = 8'hFD;
		16'hC60: out_word = 8'hCB;
		16'hC61: out_word = 8'h02;
		16'hC62: out_word = 8'h46;
		16'hC63: out_word = 8'hC2;
		16'hC64: out_word = 8'h02;
		16'hC65: out_word = 8'h0D;
		16'hC66: out_word = 8'hFD;
		16'hC67: out_word = 8'hBE;
		16'hC68: out_word = 8'h31;
		16'hC69: out_word = 8'h38;
		16'hC6A: out_word = 8'h1B;
		16'hC6B: out_word = 8'hC0;
		16'hC6C: out_word = 8'hFD;
		16'hC6D: out_word = 8'hCB;
		16'hC6E: out_word = 8'h02;
		16'hC6F: out_word = 8'h66;
		16'hC70: out_word = 8'h28;
		16'hC71: out_word = 8'h16;
		16'hC72: out_word = 8'hFD;
		16'hC73: out_word = 8'h5E;
		16'hC74: out_word = 8'h2D;
		16'hC75: out_word = 8'h1D;
		16'hC76: out_word = 8'h28;
		16'hC77: out_word = 8'h5A;
		16'hC78: out_word = 8'h3E;
		16'hC79: out_word = 8'h00;
		16'hC7A: out_word = 8'hCD;
		16'hC7B: out_word = 8'h01;
		16'hC7C: out_word = 8'h16;
		16'hC7D: out_word = 8'hED;
		16'hC7E: out_word = 8'h7B;
		16'hC7F: out_word = 8'h3F;
		16'hC80: out_word = 8'h5C;
		16'hC81: out_word = 8'hFD;
		16'hC82: out_word = 8'hCB;
		16'hC83: out_word = 8'h02;
		16'hC84: out_word = 8'hA6;
		16'hC85: out_word = 8'hC9;
		16'hC86: out_word = 8'hCF;
		16'hC87: out_word = 8'h04;
		16'hC88: out_word = 8'hFD;
		16'hC89: out_word = 8'h35;
		16'hC8A: out_word = 8'h52;
		16'hC8B: out_word = 8'h20;
		16'hC8C: out_word = 8'h45;
		16'hC8D: out_word = 8'h3E;
		16'hC8E: out_word = 8'h18;
		16'hC8F: out_word = 8'h90;
		16'hC90: out_word = 8'h32;
		16'hC91: out_word = 8'h8C;
		16'hC92: out_word = 8'h5C;
		16'hC93: out_word = 8'h2A;
		16'hC94: out_word = 8'h8F;
		16'hC95: out_word = 8'h5C;
		16'hC96: out_word = 8'hE5;
		16'hC97: out_word = 8'h3A;
		16'hC98: out_word = 8'h91;
		16'hC99: out_word = 8'h5C;
		16'hC9A: out_word = 8'hF5;
		16'hC9B: out_word = 8'h3E;
		16'hC9C: out_word = 8'hFD;
		16'hC9D: out_word = 8'hCD;
		16'hC9E: out_word = 8'h01;
		16'hC9F: out_word = 8'h16;
		16'hCA0: out_word = 8'hAF;
		16'hCA1: out_word = 8'h11;
		16'hCA2: out_word = 8'hF8;
		16'hCA3: out_word = 8'h0C;
		16'hCA4: out_word = 8'hCD;
		16'hCA5: out_word = 8'h0A;
		16'hCA6: out_word = 8'h0C;
		16'hCA7: out_word = 8'hFD;
		16'hCA8: out_word = 8'hCB;
		16'hCA9: out_word = 8'h02;
		16'hCAA: out_word = 8'hEE;
		16'hCAB: out_word = 8'h21;
		16'hCAC: out_word = 8'h3B;
		16'hCAD: out_word = 8'h5C;
		16'hCAE: out_word = 8'hCB;
		16'hCAF: out_word = 8'hDE;
		16'hCB0: out_word = 8'hCB;
		16'hCB1: out_word = 8'hAE;
		16'hCB2: out_word = 8'hD9;
		16'hCB3: out_word = 8'hCD;
		16'hCB4: out_word = 8'hD4;
		16'hCB5: out_word = 8'h15;
		16'hCB6: out_word = 8'hD9;
		16'hCB7: out_word = 8'hFE;
		16'hCB8: out_word = 8'h20;
		16'hCB9: out_word = 8'h28;
		16'hCBA: out_word = 8'h45;
		16'hCBB: out_word = 8'hFE;
		16'hCBC: out_word = 8'hE2;
		16'hCBD: out_word = 8'h28;
		16'hCBE: out_word = 8'h41;
		16'hCBF: out_word = 8'hF6;
		16'hCC0: out_word = 8'h20;
		16'hCC1: out_word = 8'hFE;
		16'hCC2: out_word = 8'h6E;
		16'hCC3: out_word = 8'h28;
		16'hCC4: out_word = 8'h3B;
		16'hCC5: out_word = 8'h3E;
		16'hCC6: out_word = 8'hFE;
		16'hCC7: out_word = 8'hCD;
		16'hCC8: out_word = 8'h01;
		16'hCC9: out_word = 8'h16;
		16'hCCA: out_word = 8'hF1;
		16'hCCB: out_word = 8'h32;
		16'hCCC: out_word = 8'h91;
		16'hCCD: out_word = 8'h5C;
		16'hCCE: out_word = 8'hE1;
		16'hCCF: out_word = 8'h22;
		16'hCD0: out_word = 8'h8F;
		16'hCD1: out_word = 8'h5C;
		16'hCD2: out_word = 8'hCD;
		16'hCD3: out_word = 8'hFE;
		16'hCD4: out_word = 8'h0D;
		16'hCD5: out_word = 8'hFD;
		16'hCD6: out_word = 8'h46;
		16'hCD7: out_word = 8'h31;
		16'hCD8: out_word = 8'h04;
		16'hCD9: out_word = 8'h0E;
		16'hCDA: out_word = 8'h21;
		16'hCDB: out_word = 8'hC5;
		16'hCDC: out_word = 8'hCD;
		16'hCDD: out_word = 8'h9B;
		16'hCDE: out_word = 8'h0E;
		16'hCDF: out_word = 8'h7C;
		16'hCE0: out_word = 8'h0F;
		16'hCE1: out_word = 8'h0F;
		16'hCE2: out_word = 8'h0F;
		16'hCE3: out_word = 8'hE6;
		16'hCE4: out_word = 8'h03;
		16'hCE5: out_word = 8'hF6;
		16'hCE6: out_word = 8'h58;
		16'hCE7: out_word = 8'h67;
		16'hCE8: out_word = 8'h11;
		16'hCE9: out_word = 8'hE0;
		16'hCEA: out_word = 8'h5A;
		16'hCEB: out_word = 8'h1A;
		16'hCEC: out_word = 8'h4E;
		16'hCED: out_word = 8'h06;
		16'hCEE: out_word = 8'h20;
		16'hCEF: out_word = 8'hEB;
		16'hCF0: out_word = 8'h12;
		16'hCF1: out_word = 8'h71;
		16'hCF2: out_word = 8'h13;
		16'hCF3: out_word = 8'h23;
		16'hCF4: out_word = 8'h10;
		16'hCF5: out_word = 8'hFA;
		16'hCF6: out_word = 8'hC1;
		16'hCF7: out_word = 8'hC9;
		16'hCF8: out_word = 8'h80;
		16'hCF9: out_word = 8'h73;
		16'hCFA: out_word = 8'h63;
		16'hCFB: out_word = 8'h72;
		16'hCFC: out_word = 8'h6F;
		16'hCFD: out_word = 8'h6C;
		16'hCFE: out_word = 8'h6C;
		16'hCFF: out_word = 8'hBF;
		16'hD00: out_word = 8'hCF;
		16'hD01: out_word = 8'h0C;
		16'hD02: out_word = 8'hFE;
		16'hD03: out_word = 8'h02;
		16'hD04: out_word = 8'h38;
		16'hD05: out_word = 8'h80;
		16'hD06: out_word = 8'hFD;
		16'hD07: out_word = 8'h86;
		16'hD08: out_word = 8'h31;
		16'hD09: out_word = 8'hD6;
		16'hD0A: out_word = 8'h19;
		16'hD0B: out_word = 8'hD0;
		16'hD0C: out_word = 8'hED;
		16'hD0D: out_word = 8'h44;
		16'hD0E: out_word = 8'hC5;
		16'hD0F: out_word = 8'h47;
		16'hD10: out_word = 8'h2A;
		16'hD11: out_word = 8'h8F;
		16'hD12: out_word = 8'h5C;
		16'hD13: out_word = 8'hE5;
		16'hD14: out_word = 8'h2A;
		16'hD15: out_word = 8'h91;
		16'hD16: out_word = 8'h5C;
		16'hD17: out_word = 8'hE5;
		16'hD18: out_word = 8'hCD;
		16'hD19: out_word = 8'h4D;
		16'hD1A: out_word = 8'h0D;
		16'hD1B: out_word = 8'h78;
		16'hD1C: out_word = 8'hF5;
		16'hD1D: out_word = 8'h21;
		16'hD1E: out_word = 8'h6B;
		16'hD1F: out_word = 8'h5C;
		16'hD20: out_word = 8'h46;
		16'hD21: out_word = 8'h78;
		16'hD22: out_word = 8'h3C;
		16'hD23: out_word = 8'h77;
		16'hD24: out_word = 8'h21;
		16'hD25: out_word = 8'h89;
		16'hD26: out_word = 8'h5C;
		16'hD27: out_word = 8'hBE;
		16'hD28: out_word = 8'h38;
		16'hD29: out_word = 8'h03;
		16'hD2A: out_word = 8'h34;
		16'hD2B: out_word = 8'h06;
		16'hD2C: out_word = 8'h18;
		16'hD2D: out_word = 8'hCD;
		16'hD2E: out_word = 8'h00;
		16'hD2F: out_word = 8'h0E;
		16'hD30: out_word = 8'hF1;
		16'hD31: out_word = 8'h3D;
		16'hD32: out_word = 8'h20;
		16'hD33: out_word = 8'hE8;
		16'hD34: out_word = 8'hE1;
		16'hD35: out_word = 8'hFD;
		16'hD36: out_word = 8'h75;
		16'hD37: out_word = 8'h57;
		16'hD38: out_word = 8'hE1;
		16'hD39: out_word = 8'h22;
		16'hD3A: out_word = 8'h8F;
		16'hD3B: out_word = 8'h5C;
		16'hD3C: out_word = 8'hED;
		16'hD3D: out_word = 8'h4B;
		16'hD3E: out_word = 8'h88;
		16'hD3F: out_word = 8'h5C;
		16'hD40: out_word = 8'hFD;
		16'hD41: out_word = 8'hCB;
		16'hD42: out_word = 8'h02;
		16'hD43: out_word = 8'h86;
		16'hD44: out_word = 8'hCD;
		16'hD45: out_word = 8'hD9;
		16'hD46: out_word = 8'h0D;
		16'hD47: out_word = 8'hFD;
		16'hD48: out_word = 8'hCB;
		16'hD49: out_word = 8'h02;
		16'hD4A: out_word = 8'hC6;
		16'hD4B: out_word = 8'hC1;
		16'hD4C: out_word = 8'hC9;
		16'hD4D: out_word = 8'hAF;
		16'hD4E: out_word = 8'h2A;
		16'hD4F: out_word = 8'h8D;
		16'hD50: out_word = 8'h5C;
		16'hD51: out_word = 8'hFD;
		16'hD52: out_word = 8'hCB;
		16'hD53: out_word = 8'h02;
		16'hD54: out_word = 8'h46;
		16'hD55: out_word = 8'h28;
		16'hD56: out_word = 8'h04;
		16'hD57: out_word = 8'h67;
		16'hD58: out_word = 8'hFD;
		16'hD59: out_word = 8'h6E;
		16'hD5A: out_word = 8'h0E;
		16'hD5B: out_word = 8'h22;
		16'hD5C: out_word = 8'h8F;
		16'hD5D: out_word = 8'h5C;
		16'hD5E: out_word = 8'h21;
		16'hD5F: out_word = 8'h91;
		16'hD60: out_word = 8'h5C;
		16'hD61: out_word = 8'h20;
		16'hD62: out_word = 8'h02;
		16'hD63: out_word = 8'h7E;
		16'hD64: out_word = 8'h0F;
		16'hD65: out_word = 8'hAE;
		16'hD66: out_word = 8'hE6;
		16'hD67: out_word = 8'h55;
		16'hD68: out_word = 8'hAE;
		16'hD69: out_word = 8'h77;
		16'hD6A: out_word = 8'hC9;
		16'hD6B: out_word = 8'hCD;
		16'hD6C: out_word = 8'hAF;
		16'hD6D: out_word = 8'h0D;
		16'hD6E: out_word = 8'h21;
		16'hD6F: out_word = 8'h3C;
		16'hD70: out_word = 8'h5C;
		16'hD71: out_word = 8'hCB;
		16'hD72: out_word = 8'hAE;
		16'hD73: out_word = 8'hCB;
		16'hD74: out_word = 8'hC6;
		16'hD75: out_word = 8'hCD;
		16'hD76: out_word = 8'h4D;
		16'hD77: out_word = 8'h0D;
		16'hD78: out_word = 8'hFD;
		16'hD79: out_word = 8'h46;
		16'hD7A: out_word = 8'h31;
		16'hD7B: out_word = 8'hCD;
		16'hD7C: out_word = 8'h44;
		16'hD7D: out_word = 8'h0E;
		16'hD7E: out_word = 8'h21;
		16'hD7F: out_word = 8'hC0;
		16'hD80: out_word = 8'h5A;
		16'hD81: out_word = 8'h3A;
		16'hD82: out_word = 8'h8D;
		16'hD83: out_word = 8'h5C;
		16'hD84: out_word = 8'h05;
		16'hD85: out_word = 8'h18;
		16'hD86: out_word = 8'h07;
		16'hD87: out_word = 8'h0E;
		16'hD88: out_word = 8'h20;
		16'hD89: out_word = 8'h2B;
		16'hD8A: out_word = 8'h77;
		16'hD8B: out_word = 8'h0D;
		16'hD8C: out_word = 8'h20;
		16'hD8D: out_word = 8'hFB;
		16'hD8E: out_word = 8'h10;
		16'hD8F: out_word = 8'hF7;
		16'hD90: out_word = 8'hFD;
		16'hD91: out_word = 8'h36;
		16'hD92: out_word = 8'h31;
		16'hD93: out_word = 8'h02;
		16'hD94: out_word = 8'h3E;
		16'hD95: out_word = 8'hFD;
		16'hD96: out_word = 8'hCD;
		16'hD97: out_word = 8'h01;
		16'hD98: out_word = 8'h16;
		16'hD99: out_word = 8'h2A;
		16'hD9A: out_word = 8'h51;
		16'hD9B: out_word = 8'h5C;
		16'hD9C: out_word = 8'h11;
		16'hD9D: out_word = 8'hF4;
		16'hD9E: out_word = 8'h09;
		16'hD9F: out_word = 8'hA7;
		16'hDA0: out_word = 8'h73;
		16'hDA1: out_word = 8'h23;
		16'hDA2: out_word = 8'h72;
		16'hDA3: out_word = 8'h23;
		16'hDA4: out_word = 8'h11;
		16'hDA5: out_word = 8'hA8;
		16'hDA6: out_word = 8'h10;
		16'hDA7: out_word = 8'h3F;
		16'hDA8: out_word = 8'h38;
		16'hDA9: out_word = 8'hF6;
		16'hDAA: out_word = 8'h01;
		16'hDAB: out_word = 8'h21;
		16'hDAC: out_word = 8'h17;
		16'hDAD: out_word = 8'h18;
		16'hDAE: out_word = 8'h2A;
		16'hDAF: out_word = 8'h21;
		16'hDB0: out_word = 8'h00;
		16'hDB1: out_word = 8'h00;
		16'hDB2: out_word = 8'h22;
		16'hDB3: out_word = 8'h7D;
		16'hDB4: out_word = 8'h5C;
		16'hDB5: out_word = 8'hFD;
		16'hDB6: out_word = 8'hCB;
		16'hDB7: out_word = 8'h30;
		16'hDB8: out_word = 8'h86;
		16'hDB9: out_word = 8'hCD;
		16'hDBA: out_word = 8'h94;
		16'hDBB: out_word = 8'h0D;
		16'hDBC: out_word = 8'h3E;
		16'hDBD: out_word = 8'hFE;
		16'hDBE: out_word = 8'hCD;
		16'hDBF: out_word = 8'h01;
		16'hDC0: out_word = 8'h16;
		16'hDC1: out_word = 8'hCD;
		16'hDC2: out_word = 8'h4D;
		16'hDC3: out_word = 8'h0D;
		16'hDC4: out_word = 8'h06;
		16'hDC5: out_word = 8'h18;
		16'hDC6: out_word = 8'hCD;
		16'hDC7: out_word = 8'h44;
		16'hDC8: out_word = 8'h0E;
		16'hDC9: out_word = 8'h2A;
		16'hDCA: out_word = 8'h51;
		16'hDCB: out_word = 8'h5C;
		16'hDCC: out_word = 8'h11;
		16'hDCD: out_word = 8'hF4;
		16'hDCE: out_word = 8'h09;
		16'hDCF: out_word = 8'h73;
		16'hDD0: out_word = 8'h23;
		16'hDD1: out_word = 8'h72;
		16'hDD2: out_word = 8'hFD;
		16'hDD3: out_word = 8'h36;
		16'hDD4: out_word = 8'h52;
		16'hDD5: out_word = 8'h01;
		16'hDD6: out_word = 8'h01;
		16'hDD7: out_word = 8'h21;
		16'hDD8: out_word = 8'h18;
		16'hDD9: out_word = 8'h21;
		16'hDDA: out_word = 8'h00;
		16'hDDB: out_word = 8'h5B;
		16'hDDC: out_word = 8'hFD;
		16'hDDD: out_word = 8'hCB;
		16'hDDE: out_word = 8'h01;
		16'hDDF: out_word = 8'h4E;
		16'hDE0: out_word = 8'h20;
		16'hDE1: out_word = 8'h12;
		16'hDE2: out_word = 8'h78;
		16'hDE3: out_word = 8'hFD;
		16'hDE4: out_word = 8'hCB;
		16'hDE5: out_word = 8'h02;
		16'hDE6: out_word = 8'h46;
		16'hDE7: out_word = 8'h28;
		16'hDE8: out_word = 8'h05;
		16'hDE9: out_word = 8'hFD;
		16'hDEA: out_word = 8'h86;
		16'hDEB: out_word = 8'h31;
		16'hDEC: out_word = 8'hD6;
		16'hDED: out_word = 8'h18;
		16'hDEE: out_word = 8'hC5;
		16'hDEF: out_word = 8'h47;
		16'hDF0: out_word = 8'hCD;
		16'hDF1: out_word = 8'h9B;
		16'hDF2: out_word = 8'h0E;
		16'hDF3: out_word = 8'hC1;
		16'hDF4: out_word = 8'h3E;
		16'hDF5: out_word = 8'h21;
		16'hDF6: out_word = 8'h91;
		16'hDF7: out_word = 8'h5F;
		16'hDF8: out_word = 8'h16;
		16'hDF9: out_word = 8'h00;
		16'hDFA: out_word = 8'h19;
		16'hDFB: out_word = 8'hC3;
		16'hDFC: out_word = 8'hDC;
		16'hDFD: out_word = 8'h0A;
		16'hDFE: out_word = 8'h06;
		16'hDFF: out_word = 8'h17;
		16'hE00: out_word = 8'hCD;
		16'hE01: out_word = 8'h9B;
		16'hE02: out_word = 8'h0E;
		16'hE03: out_word = 8'h0E;
		16'hE04: out_word = 8'h08;
		16'hE05: out_word = 8'hC5;
		16'hE06: out_word = 8'hE5;
		16'hE07: out_word = 8'h78;
		16'hE08: out_word = 8'hE6;
		16'hE09: out_word = 8'h07;
		16'hE0A: out_word = 8'h78;
		16'hE0B: out_word = 8'h20;
		16'hE0C: out_word = 8'h0C;
		16'hE0D: out_word = 8'hEB;
		16'hE0E: out_word = 8'h21;
		16'hE0F: out_word = 8'hE0;
		16'hE10: out_word = 8'hF8;
		16'hE11: out_word = 8'h19;
		16'hE12: out_word = 8'hEB;
		16'hE13: out_word = 8'h01;
		16'hE14: out_word = 8'h20;
		16'hE15: out_word = 8'h00;
		16'hE16: out_word = 8'h3D;
		16'hE17: out_word = 8'hED;
		16'hE18: out_word = 8'hB0;
		16'hE19: out_word = 8'hEB;
		16'hE1A: out_word = 8'h21;
		16'hE1B: out_word = 8'hE0;
		16'hE1C: out_word = 8'hFF;
		16'hE1D: out_word = 8'h19;
		16'hE1E: out_word = 8'hEB;
		16'hE1F: out_word = 8'h47;
		16'hE20: out_word = 8'hE6;
		16'hE21: out_word = 8'h07;
		16'hE22: out_word = 8'h0F;
		16'hE23: out_word = 8'h0F;
		16'hE24: out_word = 8'h0F;
		16'hE25: out_word = 8'h4F;
		16'hE26: out_word = 8'h78;
		16'hE27: out_word = 8'h06;
		16'hE28: out_word = 8'h00;
		16'hE29: out_word = 8'hED;
		16'hE2A: out_word = 8'hB0;
		16'hE2B: out_word = 8'h06;
		16'hE2C: out_word = 8'h07;
		16'hE2D: out_word = 8'h09;
		16'hE2E: out_word = 8'hE6;
		16'hE2F: out_word = 8'hF8;
		16'hE30: out_word = 8'h20;
		16'hE31: out_word = 8'hDB;
		16'hE32: out_word = 8'hE1;
		16'hE33: out_word = 8'h24;
		16'hE34: out_word = 8'hC1;
		16'hE35: out_word = 8'h0D;
		16'hE36: out_word = 8'h20;
		16'hE37: out_word = 8'hCD;
		16'hE38: out_word = 8'hCD;
		16'hE39: out_word = 8'h88;
		16'hE3A: out_word = 8'h0E;
		16'hE3B: out_word = 8'h21;
		16'hE3C: out_word = 8'hE0;
		16'hE3D: out_word = 8'hFF;
		16'hE3E: out_word = 8'h19;
		16'hE3F: out_word = 8'hEB;
		16'hE40: out_word = 8'hED;
		16'hE41: out_word = 8'hB0;
		16'hE42: out_word = 8'h06;
		16'hE43: out_word = 8'h01;
		16'hE44: out_word = 8'hC5;
		16'hE45: out_word = 8'hCD;
		16'hE46: out_word = 8'h9B;
		16'hE47: out_word = 8'h0E;
		16'hE48: out_word = 8'h0E;
		16'hE49: out_word = 8'h08;
		16'hE4A: out_word = 8'hC5;
		16'hE4B: out_word = 8'hE5;
		16'hE4C: out_word = 8'h78;
		16'hE4D: out_word = 8'hE6;
		16'hE4E: out_word = 8'h07;
		16'hE4F: out_word = 8'h0F;
		16'hE50: out_word = 8'h0F;
		16'hE51: out_word = 8'h0F;
		16'hE52: out_word = 8'h4F;
		16'hE53: out_word = 8'h78;
		16'hE54: out_word = 8'h06;
		16'hE55: out_word = 8'h00;
		16'hE56: out_word = 8'h0D;
		16'hE57: out_word = 8'h54;
		16'hE58: out_word = 8'h5D;
		16'hE59: out_word = 8'h36;
		16'hE5A: out_word = 8'h00;
		16'hE5B: out_word = 8'h13;
		16'hE5C: out_word = 8'hED;
		16'hE5D: out_word = 8'hB0;
		16'hE5E: out_word = 8'h11;
		16'hE5F: out_word = 8'h01;
		16'hE60: out_word = 8'h07;
		16'hE61: out_word = 8'h19;
		16'hE62: out_word = 8'h3D;
		16'hE63: out_word = 8'hE6;
		16'hE64: out_word = 8'hF8;
		16'hE65: out_word = 8'h47;
		16'hE66: out_word = 8'h20;
		16'hE67: out_word = 8'hE5;
		16'hE68: out_word = 8'hE1;
		16'hE69: out_word = 8'h24;
		16'hE6A: out_word = 8'hC1;
		16'hE6B: out_word = 8'h0D;
		16'hE6C: out_word = 8'h20;
		16'hE6D: out_word = 8'hDC;
		16'hE6E: out_word = 8'hCD;
		16'hE6F: out_word = 8'h88;
		16'hE70: out_word = 8'h0E;
		16'hE71: out_word = 8'h62;
		16'hE72: out_word = 8'h6B;
		16'hE73: out_word = 8'h13;
		16'hE74: out_word = 8'h3A;
		16'hE75: out_word = 8'h8D;
		16'hE76: out_word = 8'h5C;
		16'hE77: out_word = 8'hFD;
		16'hE78: out_word = 8'hCB;
		16'hE79: out_word = 8'h02;
		16'hE7A: out_word = 8'h46;
		16'hE7B: out_word = 8'h28;
		16'hE7C: out_word = 8'h03;
		16'hE7D: out_word = 8'h3A;
		16'hE7E: out_word = 8'h48;
		16'hE7F: out_word = 8'h5C;
		16'hE80: out_word = 8'h77;
		16'hE81: out_word = 8'h0B;
		16'hE82: out_word = 8'hED;
		16'hE83: out_word = 8'hB0;
		16'hE84: out_word = 8'hC1;
		16'hE85: out_word = 8'h0E;
		16'hE86: out_word = 8'h21;
		16'hE87: out_word = 8'hC9;
		16'hE88: out_word = 8'h7C;
		16'hE89: out_word = 8'h0F;
		16'hE8A: out_word = 8'h0F;
		16'hE8B: out_word = 8'h0F;
		16'hE8C: out_word = 8'h3D;
		16'hE8D: out_word = 8'hF6;
		16'hE8E: out_word = 8'h50;
		16'hE8F: out_word = 8'h67;
		16'hE90: out_word = 8'hEB;
		16'hE91: out_word = 8'h61;
		16'hE92: out_word = 8'h68;
		16'hE93: out_word = 8'h29;
		16'hE94: out_word = 8'h29;
		16'hE95: out_word = 8'h29;
		16'hE96: out_word = 8'h29;
		16'hE97: out_word = 8'h29;
		16'hE98: out_word = 8'h44;
		16'hE99: out_word = 8'h4D;
		16'hE9A: out_word = 8'hC9;
		16'hE9B: out_word = 8'h3E;
		16'hE9C: out_word = 8'h18;
		16'hE9D: out_word = 8'h90;
		16'hE9E: out_word = 8'h57;
		16'hE9F: out_word = 8'h0F;
		16'hEA0: out_word = 8'h0F;
		16'hEA1: out_word = 8'h0F;
		16'hEA2: out_word = 8'hE6;
		16'hEA3: out_word = 8'hE0;
		16'hEA4: out_word = 8'h6F;
		16'hEA5: out_word = 8'h7A;
		16'hEA6: out_word = 8'hE6;
		16'hEA7: out_word = 8'h18;
		16'hEA8: out_word = 8'hF6;
		16'hEA9: out_word = 8'h40;
		16'hEAA: out_word = 8'h67;
		16'hEAB: out_word = 8'hC9;
		16'hEAC: out_word = 8'hF3;
		16'hEAD: out_word = 8'h06;
		16'hEAE: out_word = 8'hB0;
		16'hEAF: out_word = 8'h21;
		16'hEB0: out_word = 8'h00;
		16'hEB1: out_word = 8'h40;
		16'hEB2: out_word = 8'hE5;
		16'hEB3: out_word = 8'hC5;
		16'hEB4: out_word = 8'hCD;
		16'hEB5: out_word = 8'hF4;
		16'hEB6: out_word = 8'h0E;
		16'hEB7: out_word = 8'hC1;
		16'hEB8: out_word = 8'hE1;
		16'hEB9: out_word = 8'h24;
		16'hEBA: out_word = 8'h7C;
		16'hEBB: out_word = 8'hE6;
		16'hEBC: out_word = 8'h07;
		16'hEBD: out_word = 8'h20;
		16'hEBE: out_word = 8'h0A;
		16'hEBF: out_word = 8'h7D;
		16'hEC0: out_word = 8'hC6;
		16'hEC1: out_word = 8'h20;
		16'hEC2: out_word = 8'h6F;
		16'hEC3: out_word = 8'h3F;
		16'hEC4: out_word = 8'h9F;
		16'hEC5: out_word = 8'hE6;
		16'hEC6: out_word = 8'hF8;
		16'hEC7: out_word = 8'h84;
		16'hEC8: out_word = 8'h67;
		16'hEC9: out_word = 8'h10;
		16'hECA: out_word = 8'hE7;
		16'hECB: out_word = 8'h18;
		16'hECC: out_word = 8'h0D;
		16'hECD: out_word = 8'hF3;
		16'hECE: out_word = 8'h21;
		16'hECF: out_word = 8'h00;
		16'hED0: out_word = 8'h5B;
		16'hED1: out_word = 8'h06;
		16'hED2: out_word = 8'h08;
		16'hED3: out_word = 8'hC5;
		16'hED4: out_word = 8'hCD;
		16'hED5: out_word = 8'hF4;
		16'hED6: out_word = 8'h0E;
		16'hED7: out_word = 8'hC1;
		16'hED8: out_word = 8'h10;
		16'hED9: out_word = 8'hF9;
		16'hEDA: out_word = 8'h3E;
		16'hEDB: out_word = 8'h04;
		16'hEDC: out_word = 8'hD3;
		16'hEDD: out_word = 8'hFB;
		16'hEDE: out_word = 8'hFB;
		16'hEDF: out_word = 8'h21;
		16'hEE0: out_word = 8'h00;
		16'hEE1: out_word = 8'h5B;
		16'hEE2: out_word = 8'hFD;
		16'hEE3: out_word = 8'h75;
		16'hEE4: out_word = 8'h46;
		16'hEE5: out_word = 8'hAF;
		16'hEE6: out_word = 8'h47;
		16'hEE7: out_word = 8'h77;
		16'hEE8: out_word = 8'h23;
		16'hEE9: out_word = 8'h10;
		16'hEEA: out_word = 8'hFC;
		16'hEEB: out_word = 8'hFD;
		16'hEEC: out_word = 8'hCB;
		16'hEED: out_word = 8'h30;
		16'hEEE: out_word = 8'h8E;
		16'hEEF: out_word = 8'h0E;
		16'hEF0: out_word = 8'h21;
		16'hEF1: out_word = 8'hC3;
		16'hEF2: out_word = 8'hD9;
		16'hEF3: out_word = 8'h0D;
		16'hEF4: out_word = 8'h78;
		16'hEF5: out_word = 8'hFE;
		16'hEF6: out_word = 8'h03;
		16'hEF7: out_word = 8'h9F;
		16'hEF8: out_word = 8'hE6;
		16'hEF9: out_word = 8'h02;
		16'hEFA: out_word = 8'hD3;
		16'hEFB: out_word = 8'hFB;
		16'hEFC: out_word = 8'h57;
		16'hEFD: out_word = 8'hCD;
		16'hEFE: out_word = 8'h54;
		16'hEFF: out_word = 8'h1F;
		16'hF00: out_word = 8'h38;
		16'hF01: out_word = 8'h0A;
		16'hF02: out_word = 8'h3E;
		16'hF03: out_word = 8'h04;
		16'hF04: out_word = 8'hD3;
		16'hF05: out_word = 8'hFB;
		16'hF06: out_word = 8'hFB;
		16'hF07: out_word = 8'hCD;
		16'hF08: out_word = 8'hDF;
		16'hF09: out_word = 8'h0E;
		16'hF0A: out_word = 8'hCF;
		16'hF0B: out_word = 8'h0C;
		16'hF0C: out_word = 8'hDB;
		16'hF0D: out_word = 8'hFB;
		16'hF0E: out_word = 8'h87;
		16'hF0F: out_word = 8'hF8;
		16'hF10: out_word = 8'h30;
		16'hF11: out_word = 8'hEB;
		16'hF12: out_word = 8'h0E;
		16'hF13: out_word = 8'h20;
		16'hF14: out_word = 8'h5E;
		16'hF15: out_word = 8'h23;
		16'hF16: out_word = 8'h06;
		16'hF17: out_word = 8'h08;
		16'hF18: out_word = 8'hCB;
		16'hF19: out_word = 8'h12;
		16'hF1A: out_word = 8'hCB;
		16'hF1B: out_word = 8'h13;
		16'hF1C: out_word = 8'hCB;
		16'hF1D: out_word = 8'h1A;
		16'hF1E: out_word = 8'hDB;
		16'hF1F: out_word = 8'hFB;
		16'hF20: out_word = 8'h1F;
		16'hF21: out_word = 8'h30;
		16'hF22: out_word = 8'hFB;
		16'hF23: out_word = 8'h7A;
		16'hF24: out_word = 8'hD3;
		16'hF25: out_word = 8'hFB;
		16'hF26: out_word = 8'h10;
		16'hF27: out_word = 8'hF0;
		16'hF28: out_word = 8'h0D;
		16'hF29: out_word = 8'h20;
		16'hF2A: out_word = 8'hE9;
		16'hF2B: out_word = 8'hC9;
		16'hF2C: out_word = 8'h2A;
		16'hF2D: out_word = 8'h3D;
		16'hF2E: out_word = 8'h5C;
		16'hF2F: out_word = 8'hE5;
		16'hF30: out_word = 8'h21;
		16'hF31: out_word = 8'h7F;
		16'hF32: out_word = 8'h10;
		16'hF33: out_word = 8'hE5;
		16'hF34: out_word = 8'hED;
		16'hF35: out_word = 8'h73;
		16'hF36: out_word = 8'h3D;
		16'hF37: out_word = 8'h5C;
		16'hF38: out_word = 8'hCD;
		16'hF39: out_word = 8'hD4;
		16'hF3A: out_word = 8'h15;
		16'hF3B: out_word = 8'hF5;
		16'hF3C: out_word = 8'h16;
		16'hF3D: out_word = 8'h00;
		16'hF3E: out_word = 8'hFD;
		16'hF3F: out_word = 8'h5E;
		16'hF40: out_word = 8'hFF;
		16'hF41: out_word = 8'h21;
		16'hF42: out_word = 8'hC8;
		16'hF43: out_word = 8'h00;
		16'hF44: out_word = 8'hCD;
		16'hF45: out_word = 8'hB5;
		16'hF46: out_word = 8'h03;
		16'hF47: out_word = 8'hF1;
		16'hF48: out_word = 8'h21;
		16'hF49: out_word = 8'h38;
		16'hF4A: out_word = 8'h0F;
		16'hF4B: out_word = 8'hE5;
		16'hF4C: out_word = 8'hFE;
		16'hF4D: out_word = 8'h18;
		16'hF4E: out_word = 8'h30;
		16'hF4F: out_word = 8'h31;
		16'hF50: out_word = 8'hFE;
		16'hF51: out_word = 8'h07;
		16'hF52: out_word = 8'h38;
		16'hF53: out_word = 8'h2D;
		16'hF54: out_word = 8'hFE;
		16'hF55: out_word = 8'h10;
		16'hF56: out_word = 8'h38;
		16'hF57: out_word = 8'h3A;
		16'hF58: out_word = 8'h01;
		16'hF59: out_word = 8'h02;
		16'hF5A: out_word = 8'h00;
		16'hF5B: out_word = 8'h57;
		16'hF5C: out_word = 8'hFE;
		16'hF5D: out_word = 8'h16;
		16'hF5E: out_word = 8'h38;
		16'hF5F: out_word = 8'h0C;
		16'hF60: out_word = 8'h03;
		16'hF61: out_word = 8'hFD;
		16'hF62: out_word = 8'hCB;
		16'hF63: out_word = 8'h37;
		16'hF64: out_word = 8'h7E;
		16'hF65: out_word = 8'hCA;
		16'hF66: out_word = 8'h1E;
		16'hF67: out_word = 8'h10;
		16'hF68: out_word = 8'hCD;
		16'hF69: out_word = 8'hD4;
		16'hF6A: out_word = 8'h15;
		16'hF6B: out_word = 8'h5F;
		16'hF6C: out_word = 8'hCD;
		16'hF6D: out_word = 8'hD4;
		16'hF6E: out_word = 8'h15;
		16'hF6F: out_word = 8'hD5;
		16'hF70: out_word = 8'h2A;
		16'hF71: out_word = 8'h5B;
		16'hF72: out_word = 8'h5C;
		16'hF73: out_word = 8'hFD;
		16'hF74: out_word = 8'hCB;
		16'hF75: out_word = 8'h07;
		16'hF76: out_word = 8'h86;
		16'hF77: out_word = 8'hCD;
		16'hF78: out_word = 8'h55;
		16'hF79: out_word = 8'h16;
		16'hF7A: out_word = 8'hC1;
		16'hF7B: out_word = 8'h23;
		16'hF7C: out_word = 8'h70;
		16'hF7D: out_word = 8'h23;
		16'hF7E: out_word = 8'h71;
		16'hF7F: out_word = 8'h18;
		16'hF80: out_word = 8'h0A;
		16'hF81: out_word = 8'hFD;
		16'hF82: out_word = 8'hCB;
		16'hF83: out_word = 8'h07;
		16'hF84: out_word = 8'h86;
		16'hF85: out_word = 8'h2A;
		16'hF86: out_word = 8'h5B;
		16'hF87: out_word = 8'h5C;
		16'hF88: out_word = 8'hCD;
		16'hF89: out_word = 8'h52;
		16'hF8A: out_word = 8'h16;
		16'hF8B: out_word = 8'h12;
		16'hF8C: out_word = 8'h13;
		16'hF8D: out_word = 8'hED;
		16'hF8E: out_word = 8'h53;
		16'hF8F: out_word = 8'h5B;
		16'hF90: out_word = 8'h5C;
		16'hF91: out_word = 8'hC9;
		16'hF92: out_word = 8'h5F;
		16'hF93: out_word = 8'h16;
		16'hF94: out_word = 8'h00;
		16'hF95: out_word = 8'h21;
		16'hF96: out_word = 8'h99;
		16'hF97: out_word = 8'h0F;
		16'hF98: out_word = 8'h19;
		16'hF99: out_word = 8'h5E;
		16'hF9A: out_word = 8'h19;
		16'hF9B: out_word = 8'hE5;
		16'hF9C: out_word = 8'h2A;
		16'hF9D: out_word = 8'h5B;
		16'hF9E: out_word = 8'h5C;
		16'hF9F: out_word = 8'hC9;
		16'hFA0: out_word = 8'h09;
		16'hFA1: out_word = 8'h66;
		16'hFA2: out_word = 8'h6A;
		16'hFA3: out_word = 8'h50;
		16'hFA4: out_word = 8'hB5;
		16'hFA5: out_word = 8'h70;
		16'hFA6: out_word = 8'h7E;
		16'hFA7: out_word = 8'hCF;
		16'hFA8: out_word = 8'hD4;
		16'hFA9: out_word = 8'h2A;
		16'hFAA: out_word = 8'h49;
		16'hFAB: out_word = 8'h5C;
		16'hFAC: out_word = 8'hFD;
		16'hFAD: out_word = 8'hCB;
		16'hFAE: out_word = 8'h37;
		16'hFAF: out_word = 8'h6E;
		16'hFB0: out_word = 8'hC2;
		16'hFB1: out_word = 8'h97;
		16'hFB2: out_word = 8'h10;
		16'hFB3: out_word = 8'hCD;
		16'hFB4: out_word = 8'h6E;
		16'hFB5: out_word = 8'h19;
		16'hFB6: out_word = 8'hCD;
		16'hFB7: out_word = 8'h95;
		16'hFB8: out_word = 8'h16;
		16'hFB9: out_word = 8'h7A;
		16'hFBA: out_word = 8'hB3;
		16'hFBB: out_word = 8'hCA;
		16'hFBC: out_word = 8'h97;
		16'hFBD: out_word = 8'h10;
		16'hFBE: out_word = 8'hE5;
		16'hFBF: out_word = 8'h23;
		16'hFC0: out_word = 8'h4E;
		16'hFC1: out_word = 8'h23;
		16'hFC2: out_word = 8'h46;
		16'hFC3: out_word = 8'h21;
		16'hFC4: out_word = 8'h0A;
		16'hFC5: out_word = 8'h00;
		16'hFC6: out_word = 8'h09;
		16'hFC7: out_word = 8'h44;
		16'hFC8: out_word = 8'h4D;
		16'hFC9: out_word = 8'hCD;
		16'hFCA: out_word = 8'h05;
		16'hFCB: out_word = 8'h1F;
		16'hFCC: out_word = 8'hCD;
		16'hFCD: out_word = 8'h97;
		16'hFCE: out_word = 8'h10;
		16'hFCF: out_word = 8'h2A;
		16'hFD0: out_word = 8'h51;
		16'hFD1: out_word = 8'h5C;
		16'hFD2: out_word = 8'hE3;
		16'hFD3: out_word = 8'hE5;
		16'hFD4: out_word = 8'h3E;
		16'hFD5: out_word = 8'hFF;
		16'hFD6: out_word = 8'hCD;
		16'hFD7: out_word = 8'h01;
		16'hFD8: out_word = 8'h16;
		16'hFD9: out_word = 8'hE1;
		16'hFDA: out_word = 8'h2B;
		16'hFDB: out_word = 8'hFD;
		16'hFDC: out_word = 8'h35;
		16'hFDD: out_word = 8'h0F;
		16'hFDE: out_word = 8'hCD;
		16'hFDF: out_word = 8'h55;
		16'hFE0: out_word = 8'h18;
		16'hFE1: out_word = 8'hFD;
		16'hFE2: out_word = 8'h34;
		16'hFE3: out_word = 8'h0F;
		16'hFE4: out_word = 8'h2A;
		16'hFE5: out_word = 8'h59;
		16'hFE6: out_word = 8'h5C;
		16'hFE7: out_word = 8'h23;
		16'hFE8: out_word = 8'h23;
		16'hFE9: out_word = 8'h23;
		16'hFEA: out_word = 8'h23;
		16'hFEB: out_word = 8'h22;
		16'hFEC: out_word = 8'h5B;
		16'hFED: out_word = 8'h5C;
		16'hFEE: out_word = 8'hE1;
		16'hFEF: out_word = 8'hCD;
		16'hFF0: out_word = 8'h15;
		16'hFF1: out_word = 8'h16;
		16'hFF2: out_word = 8'hC9;
		16'hFF3: out_word = 8'hFD;
		16'hFF4: out_word = 8'hCB;
		16'hFF5: out_word = 8'h37;
		16'hFF6: out_word = 8'h6E;
		16'hFF7: out_word = 8'h20;
		16'hFF8: out_word = 8'h08;
		16'hFF9: out_word = 8'h21;
		16'hFFA: out_word = 8'h49;
		16'hFFB: out_word = 8'h5C;
		16'hFFC: out_word = 8'hCD;
		16'hFFD: out_word = 8'h0F;
		16'hFFE: out_word = 8'h19;
		16'hFFF: out_word = 8'h18;
		16'h1000: out_word = 8'h6D;
		16'h1001: out_word = 8'hFD;
		16'h1002: out_word = 8'h36;
		16'h1003: out_word = 8'h00;
		16'h1004: out_word = 8'h10;
		16'h1005: out_word = 8'h18;
		16'h1006: out_word = 8'h1D;
		16'h1007: out_word = 8'hCD;
		16'h1008: out_word = 8'h31;
		16'h1009: out_word = 8'h10;
		16'h100A: out_word = 8'h18;
		16'h100B: out_word = 8'h05;
		16'h100C: out_word = 8'h7E;
		16'h100D: out_word = 8'hFE;
		16'h100E: out_word = 8'h0D;
		16'h100F: out_word = 8'hC8;
		16'h1010: out_word = 8'h23;
		16'h1011: out_word = 8'h22;
		16'h1012: out_word = 8'h5B;
		16'h1013: out_word = 8'h5C;
		16'h1014: out_word = 8'hC9;
		16'h1015: out_word = 8'hCD;
		16'h1016: out_word = 8'h31;
		16'h1017: out_word = 8'h10;
		16'h1018: out_word = 8'h01;
		16'h1019: out_word = 8'h01;
		16'h101A: out_word = 8'h00;
		16'h101B: out_word = 8'hC3;
		16'h101C: out_word = 8'hE8;
		16'h101D: out_word = 8'h19;
		16'h101E: out_word = 8'hCD;
		16'h101F: out_word = 8'hD4;
		16'h1020: out_word = 8'h15;
		16'h1021: out_word = 8'hCD;
		16'h1022: out_word = 8'hD4;
		16'h1023: out_word = 8'h15;
		16'h1024: out_word = 8'hE1;
		16'h1025: out_word = 8'hE1;
		16'h1026: out_word = 8'hE1;
		16'h1027: out_word = 8'h22;
		16'h1028: out_word = 8'h3D;
		16'h1029: out_word = 8'h5C;
		16'h102A: out_word = 8'hFD;
		16'h102B: out_word = 8'hCB;
		16'h102C: out_word = 8'h00;
		16'h102D: out_word = 8'h7E;
		16'h102E: out_word = 8'hC0;
		16'h102F: out_word = 8'hF9;
		16'h1030: out_word = 8'hC9;
		16'h1031: out_word = 8'h37;
		16'h1032: out_word = 8'hCD;
		16'h1033: out_word = 8'h95;
		16'h1034: out_word = 8'h11;
		16'h1035: out_word = 8'hED;
		16'h1036: out_word = 8'h52;
		16'h1037: out_word = 8'h19;
		16'h1038: out_word = 8'h23;
		16'h1039: out_word = 8'hC1;
		16'h103A: out_word = 8'hD8;
		16'h103B: out_word = 8'hC5;
		16'h103C: out_word = 8'h44;
		16'h103D: out_word = 8'h4D;
		16'h103E: out_word = 8'h62;
		16'h103F: out_word = 8'h6B;
		16'h1040: out_word = 8'h23;
		16'h1041: out_word = 8'h1A;
		16'h1042: out_word = 8'hE6;
		16'h1043: out_word = 8'hF0;
		16'h1044: out_word = 8'hFE;
		16'h1045: out_word = 8'h10;
		16'h1046: out_word = 8'h20;
		16'h1047: out_word = 8'h09;
		16'h1048: out_word = 8'h23;
		16'h1049: out_word = 8'h1A;
		16'h104A: out_word = 8'hD6;
		16'h104B: out_word = 8'h17;
		16'h104C: out_word = 8'hCE;
		16'h104D: out_word = 8'h00;
		16'h104E: out_word = 8'h20;
		16'h104F: out_word = 8'h01;
		16'h1050: out_word = 8'h23;
		16'h1051: out_word = 8'hA7;
		16'h1052: out_word = 8'hED;
		16'h1053: out_word = 8'h42;
		16'h1054: out_word = 8'h09;
		16'h1055: out_word = 8'hEB;
		16'h1056: out_word = 8'h38;
		16'h1057: out_word = 8'hE6;
		16'h1058: out_word = 8'hC9;
		16'h1059: out_word = 8'hFD;
		16'h105A: out_word = 8'hCB;
		16'h105B: out_word = 8'h37;
		16'h105C: out_word = 8'h6E;
		16'h105D: out_word = 8'hC0;
		16'h105E: out_word = 8'h2A;
		16'h105F: out_word = 8'h49;
		16'h1060: out_word = 8'h5C;
		16'h1061: out_word = 8'hCD;
		16'h1062: out_word = 8'h6E;
		16'h1063: out_word = 8'h19;
		16'h1064: out_word = 8'hEB;
		16'h1065: out_word = 8'hCD;
		16'h1066: out_word = 8'h95;
		16'h1067: out_word = 8'h16;
		16'h1068: out_word = 8'h21;
		16'h1069: out_word = 8'h4A;
		16'h106A: out_word = 8'h5C;
		16'h106B: out_word = 8'hCD;
		16'h106C: out_word = 8'h1C;
		16'h106D: out_word = 8'h19;
		16'h106E: out_word = 8'hCD;
		16'h106F: out_word = 8'h95;
		16'h1070: out_word = 8'h17;
		16'h1071: out_word = 8'h3E;
		16'h1072: out_word = 8'h00;
		16'h1073: out_word = 8'hC3;
		16'h1074: out_word = 8'h01;
		16'h1075: out_word = 8'h16;
		16'h1076: out_word = 8'hFD;
		16'h1077: out_word = 8'hCB;
		16'h1078: out_word = 8'h37;
		16'h1079: out_word = 8'h7E;
		16'h107A: out_word = 8'h28;
		16'h107B: out_word = 8'hA8;
		16'h107C: out_word = 8'hC3;
		16'h107D: out_word = 8'h81;
		16'h107E: out_word = 8'h0F;
		16'h107F: out_word = 8'hFD;
		16'h1080: out_word = 8'hCB;
		16'h1081: out_word = 8'h30;
		16'h1082: out_word = 8'h66;
		16'h1083: out_word = 8'h28;
		16'h1084: out_word = 8'hA1;
		16'h1085: out_word = 8'hFD;
		16'h1086: out_word = 8'h36;
		16'h1087: out_word = 8'h00;
		16'h1088: out_word = 8'hFF;
		16'h1089: out_word = 8'h16;
		16'h108A: out_word = 8'h00;
		16'h108B: out_word = 8'hFD;
		16'h108C: out_word = 8'h5E;
		16'h108D: out_word = 8'hFE;
		16'h108E: out_word = 8'h21;
		16'h108F: out_word = 8'h90;
		16'h1090: out_word = 8'h1A;
		16'h1091: out_word = 8'hCD;
		16'h1092: out_word = 8'hB5;
		16'h1093: out_word = 8'h03;
		16'h1094: out_word = 8'hC3;
		16'h1095: out_word = 8'h30;
		16'h1096: out_word = 8'h0F;
		16'h1097: out_word = 8'hE5;
		16'h1098: out_word = 8'hCD;
		16'h1099: out_word = 8'h90;
		16'h109A: out_word = 8'h11;
		16'h109B: out_word = 8'h2B;
		16'h109C: out_word = 8'hCD;
		16'h109D: out_word = 8'hE5;
		16'h109E: out_word = 8'h19;
		16'h109F: out_word = 8'h22;
		16'h10A0: out_word = 8'h5B;
		16'h10A1: out_word = 8'h5C;
		16'h10A2: out_word = 8'hFD;
		16'h10A3: out_word = 8'h36;
		16'h10A4: out_word = 8'h07;
		16'h10A5: out_word = 8'h00;
		16'h10A6: out_word = 8'hE1;
		16'h10A7: out_word = 8'hC9;
		16'h10A8: out_word = 8'hFD;
		16'h10A9: out_word = 8'hCB;
		16'h10AA: out_word = 8'h02;
		16'h10AB: out_word = 8'h5E;
		16'h10AC: out_word = 8'hC4;
		16'h10AD: out_word = 8'h1D;
		16'h10AE: out_word = 8'h11;
		16'h10AF: out_word = 8'hA7;
		16'h10B0: out_word = 8'hFD;
		16'h10B1: out_word = 8'hCB;
		16'h10B2: out_word = 8'h01;
		16'h10B3: out_word = 8'h6E;
		16'h10B4: out_word = 8'hC8;
		16'h10B5: out_word = 8'h3A;
		16'h10B6: out_word = 8'h08;
		16'h10B7: out_word = 8'h5C;
		16'h10B8: out_word = 8'hFD;
		16'h10B9: out_word = 8'hCB;
		16'h10BA: out_word = 8'h01;
		16'h10BB: out_word = 8'hAE;
		16'h10BC: out_word = 8'hF5;
		16'h10BD: out_word = 8'hFD;
		16'h10BE: out_word = 8'hCB;
		16'h10BF: out_word = 8'h02;
		16'h10C0: out_word = 8'h6E;
		16'h10C1: out_word = 8'hC4;
		16'h10C2: out_word = 8'h6E;
		16'h10C3: out_word = 8'h0D;
		16'h10C4: out_word = 8'hF1;
		16'h10C5: out_word = 8'hFE;
		16'h10C6: out_word = 8'h20;
		16'h10C7: out_word = 8'h30;
		16'h10C8: out_word = 8'h52;
		16'h10C9: out_word = 8'hFE;
		16'h10CA: out_word = 8'h10;
		16'h10CB: out_word = 8'h30;
		16'h10CC: out_word = 8'h2D;
		16'h10CD: out_word = 8'hFE;
		16'h10CE: out_word = 8'h06;
		16'h10CF: out_word = 8'h30;
		16'h10D0: out_word = 8'h0A;
		16'h10D1: out_word = 8'h47;
		16'h10D2: out_word = 8'hE6;
		16'h10D3: out_word = 8'h01;
		16'h10D4: out_word = 8'h4F;
		16'h10D5: out_word = 8'h78;
		16'h10D6: out_word = 8'h1F;
		16'h10D7: out_word = 8'hC6;
		16'h10D8: out_word = 8'h12;
		16'h10D9: out_word = 8'h18;
		16'h10DA: out_word = 8'h2A;
		16'h10DB: out_word = 8'h20;
		16'h10DC: out_word = 8'h09;
		16'h10DD: out_word = 8'h21;
		16'h10DE: out_word = 8'h6A;
		16'h10DF: out_word = 8'h5C;
		16'h10E0: out_word = 8'h3E;
		16'h10E1: out_word = 8'h08;
		16'h10E2: out_word = 8'hAE;
		16'h10E3: out_word = 8'h77;
		16'h10E4: out_word = 8'h18;
		16'h10E5: out_word = 8'h0E;
		16'h10E6: out_word = 8'hFE;
		16'h10E7: out_word = 8'h0E;
		16'h10E8: out_word = 8'hD8;
		16'h10E9: out_word = 8'hD6;
		16'h10EA: out_word = 8'h0D;
		16'h10EB: out_word = 8'h21;
		16'h10EC: out_word = 8'h41;
		16'h10ED: out_word = 8'h5C;
		16'h10EE: out_word = 8'hBE;
		16'h10EF: out_word = 8'h77;
		16'h10F0: out_word = 8'h20;
		16'h10F1: out_word = 8'h02;
		16'h10F2: out_word = 8'h36;
		16'h10F3: out_word = 8'h00;
		16'h10F4: out_word = 8'hFD;
		16'h10F5: out_word = 8'hCB;
		16'h10F6: out_word = 8'h02;
		16'h10F7: out_word = 8'hDE;
		16'h10F8: out_word = 8'hBF;
		16'h10F9: out_word = 8'hC9;
		16'h10FA: out_word = 8'h47;
		16'h10FB: out_word = 8'hE6;
		16'h10FC: out_word = 8'h07;
		16'h10FD: out_word = 8'h4F;
		16'h10FE: out_word = 8'h3E;
		16'h10FF: out_word = 8'h10;
		16'h1100: out_word = 8'hCB;
		16'h1101: out_word = 8'h58;
		16'h1102: out_word = 8'h20;
		16'h1103: out_word = 8'h01;
		16'h1104: out_word = 8'h3C;
		16'h1105: out_word = 8'hFD;
		16'h1106: out_word = 8'h71;
		16'h1107: out_word = 8'hD3;
		16'h1108: out_word = 8'h11;
		16'h1109: out_word = 8'h0D;
		16'h110A: out_word = 8'h11;
		16'h110B: out_word = 8'h18;
		16'h110C: out_word = 8'h06;
		16'h110D: out_word = 8'h3A;
		16'h110E: out_word = 8'h0D;
		16'h110F: out_word = 8'h5C;
		16'h1110: out_word = 8'h11;
		16'h1111: out_word = 8'hA8;
		16'h1112: out_word = 8'h10;
		16'h1113: out_word = 8'h2A;
		16'h1114: out_word = 8'h4F;
		16'h1115: out_word = 8'h5C;
		16'h1116: out_word = 8'h23;
		16'h1117: out_word = 8'h23;
		16'h1118: out_word = 8'h73;
		16'h1119: out_word = 8'h23;
		16'h111A: out_word = 8'h72;
		16'h111B: out_word = 8'h37;
		16'h111C: out_word = 8'hC9;
		16'h111D: out_word = 8'hCD;
		16'h111E: out_word = 8'h4D;
		16'h111F: out_word = 8'h0D;
		16'h1120: out_word = 8'hFD;
		16'h1121: out_word = 8'hCB;
		16'h1122: out_word = 8'h02;
		16'h1123: out_word = 8'h9E;
		16'h1124: out_word = 8'hFD;
		16'h1125: out_word = 8'hCB;
		16'h1126: out_word = 8'h02;
		16'h1127: out_word = 8'hAE;
		16'h1128: out_word = 8'h2A;
		16'h1129: out_word = 8'h8A;
		16'h112A: out_word = 8'h5C;
		16'h112B: out_word = 8'hE5;
		16'h112C: out_word = 8'h2A;
		16'h112D: out_word = 8'h3D;
		16'h112E: out_word = 8'h5C;
		16'h112F: out_word = 8'hE5;
		16'h1130: out_word = 8'h21;
		16'h1131: out_word = 8'h67;
		16'h1132: out_word = 8'h11;
		16'h1133: out_word = 8'hE5;
		16'h1134: out_word = 8'hED;
		16'h1135: out_word = 8'h73;
		16'h1136: out_word = 8'h3D;
		16'h1137: out_word = 8'h5C;
		16'h1138: out_word = 8'h2A;
		16'h1139: out_word = 8'h82;
		16'h113A: out_word = 8'h5C;
		16'h113B: out_word = 8'hE5;
		16'h113C: out_word = 8'h37;
		16'h113D: out_word = 8'hCD;
		16'h113E: out_word = 8'h95;
		16'h113F: out_word = 8'h11;
		16'h1140: out_word = 8'hEB;
		16'h1141: out_word = 8'hCD;
		16'h1142: out_word = 8'h7D;
		16'h1143: out_word = 8'h18;
		16'h1144: out_word = 8'hEB;
		16'h1145: out_word = 8'hCD;
		16'h1146: out_word = 8'hE1;
		16'h1147: out_word = 8'h18;
		16'h1148: out_word = 8'h2A;
		16'h1149: out_word = 8'h8A;
		16'h114A: out_word = 8'h5C;
		16'h114B: out_word = 8'hE3;
		16'h114C: out_word = 8'hEB;
		16'h114D: out_word = 8'hCD;
		16'h114E: out_word = 8'h4D;
		16'h114F: out_word = 8'h0D;
		16'h1150: out_word = 8'h3A;
		16'h1151: out_word = 8'h8B;
		16'h1152: out_word = 8'h5C;
		16'h1153: out_word = 8'h92;
		16'h1154: out_word = 8'h38;
		16'h1155: out_word = 8'h26;
		16'h1156: out_word = 8'h20;
		16'h1157: out_word = 8'h06;
		16'h1158: out_word = 8'h7B;
		16'h1159: out_word = 8'hFD;
		16'h115A: out_word = 8'h96;
		16'h115B: out_word = 8'h50;
		16'h115C: out_word = 8'h30;
		16'h115D: out_word = 8'h1E;
		16'h115E: out_word = 8'h3E;
		16'h115F: out_word = 8'h20;
		16'h1160: out_word = 8'hD5;
		16'h1161: out_word = 8'hCD;
		16'h1162: out_word = 8'hF4;
		16'h1163: out_word = 8'h09;
		16'h1164: out_word = 8'hD1;
		16'h1165: out_word = 8'h18;
		16'h1166: out_word = 8'hE9;
		16'h1167: out_word = 8'h16;
		16'h1168: out_word = 8'h00;
		16'h1169: out_word = 8'hFD;
		16'h116A: out_word = 8'h5E;
		16'h116B: out_word = 8'hFE;
		16'h116C: out_word = 8'h21;
		16'h116D: out_word = 8'h90;
		16'h116E: out_word = 8'h1A;
		16'h116F: out_word = 8'hCD;
		16'h1170: out_word = 8'hB5;
		16'h1171: out_word = 8'h03;
		16'h1172: out_word = 8'hFD;
		16'h1173: out_word = 8'h36;
		16'h1174: out_word = 8'h00;
		16'h1175: out_word = 8'hFF;
		16'h1176: out_word = 8'hED;
		16'h1177: out_word = 8'h5B;
		16'h1178: out_word = 8'h8A;
		16'h1179: out_word = 8'h5C;
		16'h117A: out_word = 8'h18;
		16'h117B: out_word = 8'h02;
		16'h117C: out_word = 8'hD1;
		16'h117D: out_word = 8'hE1;
		16'h117E: out_word = 8'hE1;
		16'h117F: out_word = 8'h22;
		16'h1180: out_word = 8'h3D;
		16'h1181: out_word = 8'h5C;
		16'h1182: out_word = 8'hC1;
		16'h1183: out_word = 8'hD5;
		16'h1184: out_word = 8'hCD;
		16'h1185: out_word = 8'hD9;
		16'h1186: out_word = 8'h0D;
		16'h1187: out_word = 8'hE1;
		16'h1188: out_word = 8'h22;
		16'h1189: out_word = 8'h82;
		16'h118A: out_word = 8'h5C;
		16'h118B: out_word = 8'hFD;
		16'h118C: out_word = 8'h36;
		16'h118D: out_word = 8'h26;
		16'h118E: out_word = 8'h00;
		16'h118F: out_word = 8'hC9;
		16'h1190: out_word = 8'h2A;
		16'h1191: out_word = 8'h61;
		16'h1192: out_word = 8'h5C;
		16'h1193: out_word = 8'h2B;
		16'h1194: out_word = 8'hA7;
		16'h1195: out_word = 8'hED;
		16'h1196: out_word = 8'h5B;
		16'h1197: out_word = 8'h59;
		16'h1198: out_word = 8'h5C;
		16'h1199: out_word = 8'hFD;
		16'h119A: out_word = 8'hCB;
		16'h119B: out_word = 8'h37;
		16'h119C: out_word = 8'h6E;
		16'h119D: out_word = 8'hC8;
		16'h119E: out_word = 8'hED;
		16'h119F: out_word = 8'h5B;
		16'h11A0: out_word = 8'h61;
		16'h11A1: out_word = 8'h5C;
		16'h11A2: out_word = 8'hD8;
		16'h11A3: out_word = 8'h2A;
		16'h11A4: out_word = 8'h63;
		16'h11A5: out_word = 8'h5C;
		16'h11A6: out_word = 8'hC9;
		16'h11A7: out_word = 8'h7E;
		16'h11A8: out_word = 8'hFE;
		16'h11A9: out_word = 8'h0E;
		16'h11AA: out_word = 8'h01;
		16'h11AB: out_word = 8'h06;
		16'h11AC: out_word = 8'h00;
		16'h11AD: out_word = 8'hCC;
		16'h11AE: out_word = 8'hE8;
		16'h11AF: out_word = 8'h19;
		16'h11B0: out_word = 8'h7E;
		16'h11B1: out_word = 8'h23;
		16'h11B2: out_word = 8'hFE;
		16'h11B3: out_word = 8'h0D;
		16'h11B4: out_word = 8'h20;
		16'h11B5: out_word = 8'hF1;
		16'h11B6: out_word = 8'hC9;
		16'h11B7: out_word = 8'hF3;
		16'h11B8: out_word = 8'h3E;
		16'h11B9: out_word = 8'hFF;
		16'h11BA: out_word = 8'hED;
		16'h11BB: out_word = 8'h5B;
		16'h11BC: out_word = 8'hB2;
		16'h11BD: out_word = 8'h5C;
		16'h11BE: out_word = 8'hD9;
		16'h11BF: out_word = 8'hED;
		16'h11C0: out_word = 8'h4B;
		16'h11C1: out_word = 8'hB4;
		16'h11C2: out_word = 8'h5C;
		16'h11C3: out_word = 8'hED;
		16'h11C4: out_word = 8'h5B;
		16'h11C5: out_word = 8'h38;
		16'h11C6: out_word = 8'h5C;
		16'h11C7: out_word = 8'h2A;
		16'h11C8: out_word = 8'h7B;
		16'h11C9: out_word = 8'h5C;
		16'h11CA: out_word = 8'hD9;
		16'h11CB: out_word = 8'h47;
		16'h11CC: out_word = 8'h3E;
		16'h11CD: out_word = 8'h07;
		16'h11CE: out_word = 8'hD3;
		16'h11CF: out_word = 8'hFE;
		16'h11D0: out_word = 8'h3E;
		16'h11D1: out_word = 8'h3F;
		16'h11D2: out_word = 8'hED;
		16'h11D3: out_word = 8'h47;
		16'h11D4: out_word = 8'h00;
		16'h11D5: out_word = 8'h00;
		16'h11D6: out_word = 8'h00;
		16'h11D7: out_word = 8'h00;
		16'h11D8: out_word = 8'h00;
		16'h11D9: out_word = 8'h00;
		16'h11DA: out_word = 8'h62;
		16'h11DB: out_word = 8'h6B;
		16'h11DC: out_word = 8'h36;
		16'h11DD: out_word = 8'h02;
		16'h11DE: out_word = 8'h2B;
		16'h11DF: out_word = 8'hBC;
		16'h11E0: out_word = 8'h20;
		16'h11E1: out_word = 8'hFA;
		16'h11E2: out_word = 8'hA7;
		16'h11E3: out_word = 8'hED;
		16'h11E4: out_word = 8'h52;
		16'h11E5: out_word = 8'h19;
		16'h11E6: out_word = 8'h23;
		16'h11E7: out_word = 8'h30;
		16'h11E8: out_word = 8'h06;
		16'h11E9: out_word = 8'h35;
		16'h11EA: out_word = 8'h28;
		16'h11EB: out_word = 8'h03;
		16'h11EC: out_word = 8'h35;
		16'h11ED: out_word = 8'h28;
		16'h11EE: out_word = 8'hF3;
		16'h11EF: out_word = 8'h2B;
		16'h11F0: out_word = 8'hD9;
		16'h11F1: out_word = 8'hED;
		16'h11F2: out_word = 8'h43;
		16'h11F3: out_word = 8'hB4;
		16'h11F4: out_word = 8'h5C;
		16'h11F5: out_word = 8'hED;
		16'h11F6: out_word = 8'h53;
		16'h11F7: out_word = 8'h38;
		16'h11F8: out_word = 8'h5C;
		16'h11F9: out_word = 8'h22;
		16'h11FA: out_word = 8'h7B;
		16'h11FB: out_word = 8'h5C;
		16'h11FC: out_word = 8'hD9;
		16'h11FD: out_word = 8'h04;
		16'h11FE: out_word = 8'h28;
		16'h11FF: out_word = 8'h19;
		16'h1200: out_word = 8'h22;
		16'h1201: out_word = 8'hB4;
		16'h1202: out_word = 8'h5C;
		16'h1203: out_word = 8'h11;
		16'h1204: out_word = 8'hAF;
		16'h1205: out_word = 8'h3E;
		16'h1206: out_word = 8'h01;
		16'h1207: out_word = 8'hA8;
		16'h1208: out_word = 8'h00;
		16'h1209: out_word = 8'hEB;
		16'h120A: out_word = 8'hED;
		16'h120B: out_word = 8'hB8;
		16'h120C: out_word = 8'hEB;
		16'h120D: out_word = 8'h23;
		16'h120E: out_word = 8'h22;
		16'h120F: out_word = 8'h7B;
		16'h1210: out_word = 8'h5C;
		16'h1211: out_word = 8'h2B;
		16'h1212: out_word = 8'h01;
		16'h1213: out_word = 8'h40;
		16'h1214: out_word = 8'h00;
		16'h1215: out_word = 8'hED;
		16'h1216: out_word = 8'h43;
		16'h1217: out_word = 8'h38;
		16'h1218: out_word = 8'h5C;
		16'h1219: out_word = 8'h22;
		16'h121A: out_word = 8'hB2;
		16'h121B: out_word = 8'h5C;
		16'h121C: out_word = 8'h21;
		16'h121D: out_word = 8'h00;
		16'h121E: out_word = 8'h3C;
		16'h121F: out_word = 8'h22;
		16'h1220: out_word = 8'h36;
		16'h1221: out_word = 8'h5C;
		16'h1222: out_word = 8'h2A;
		16'h1223: out_word = 8'hB2;
		16'h1224: out_word = 8'h5C;
		16'h1225: out_word = 8'h36;
		16'h1226: out_word = 8'h3E;
		16'h1227: out_word = 8'h2B;
		16'h1228: out_word = 8'hF9;
		16'h1229: out_word = 8'h2B;
		16'h122A: out_word = 8'h2B;
		16'h122B: out_word = 8'h22;
		16'h122C: out_word = 8'h3D;
		16'h122D: out_word = 8'h5C;
		16'h122E: out_word = 8'hED;
		16'h122F: out_word = 8'h56;
		16'h1230: out_word = 8'hFD;
		16'h1231: out_word = 8'h21;
		16'h1232: out_word = 8'h3A;
		16'h1233: out_word = 8'h5C;
		16'h1234: out_word = 8'hFB;
		16'h1235: out_word = 8'h21;
		16'h1236: out_word = 8'hB6;
		16'h1237: out_word = 8'h5C;
		16'h1238: out_word = 8'h22;
		16'h1239: out_word = 8'h4F;
		16'h123A: out_word = 8'h5C;
		16'h123B: out_word = 8'h11;
		16'h123C: out_word = 8'hAF;
		16'h123D: out_word = 8'h15;
		16'h123E: out_word = 8'h01;
		16'h123F: out_word = 8'h15;
		16'h1240: out_word = 8'h00;
		16'h1241: out_word = 8'hEB;
		16'h1242: out_word = 8'hED;
		16'h1243: out_word = 8'hB0;
		16'h1244: out_word = 8'hEB;
		16'h1245: out_word = 8'h2B;
		16'h1246: out_word = 8'h22;
		16'h1247: out_word = 8'h57;
		16'h1248: out_word = 8'h5C;
		16'h1249: out_word = 8'h23;
		16'h124A: out_word = 8'h22;
		16'h124B: out_word = 8'h53;
		16'h124C: out_word = 8'h5C;
		16'h124D: out_word = 8'h22;
		16'h124E: out_word = 8'h4B;
		16'h124F: out_word = 8'h5C;
		16'h1250: out_word = 8'h36;
		16'h1251: out_word = 8'h80;
		16'h1252: out_word = 8'h23;
		16'h1253: out_word = 8'h22;
		16'h1254: out_word = 8'h59;
		16'h1255: out_word = 8'h5C;
		16'h1256: out_word = 8'h36;
		16'h1257: out_word = 8'h0D;
		16'h1258: out_word = 8'h23;
		16'h1259: out_word = 8'h36;
		16'h125A: out_word = 8'h80;
		16'h125B: out_word = 8'h23;
		16'h125C: out_word = 8'h22;
		16'h125D: out_word = 8'h61;
		16'h125E: out_word = 8'h5C;
		16'h125F: out_word = 8'h22;
		16'h1260: out_word = 8'h63;
		16'h1261: out_word = 8'h5C;
		16'h1262: out_word = 8'h22;
		16'h1263: out_word = 8'h65;
		16'h1264: out_word = 8'h5C;
		16'h1265: out_word = 8'h3E;
		16'h1266: out_word = 8'h38;
		16'h1267: out_word = 8'h32;
		16'h1268: out_word = 8'h8D;
		16'h1269: out_word = 8'h5C;
		16'h126A: out_word = 8'h32;
		16'h126B: out_word = 8'h8F;
		16'h126C: out_word = 8'h5C;
		16'h126D: out_word = 8'h32;
		16'h126E: out_word = 8'h48;
		16'h126F: out_word = 8'h5C;
		16'h1270: out_word = 8'h21;
		16'h1271: out_word = 8'h23;
		16'h1272: out_word = 8'h05;
		16'h1273: out_word = 8'h22;
		16'h1274: out_word = 8'h09;
		16'h1275: out_word = 8'h5C;
		16'h1276: out_word = 8'hFD;
		16'h1277: out_word = 8'h35;
		16'h1278: out_word = 8'hC6;
		16'h1279: out_word = 8'hFD;
		16'h127A: out_word = 8'h35;
		16'h127B: out_word = 8'hCA;
		16'h127C: out_word = 8'h21;
		16'h127D: out_word = 8'hC6;
		16'h127E: out_word = 8'h15;
		16'h127F: out_word = 8'h11;
		16'h1280: out_word = 8'h10;
		16'h1281: out_word = 8'h5C;
		16'h1282: out_word = 8'h01;
		16'h1283: out_word = 8'h0E;
		16'h1284: out_word = 8'h00;
		16'h1285: out_word = 8'hED;
		16'h1286: out_word = 8'hB0;
		16'h1287: out_word = 8'hFD;
		16'h1288: out_word = 8'hCB;
		16'h1289: out_word = 8'h01;
		16'h128A: out_word = 8'hCE;
		16'h128B: out_word = 8'hCD;
		16'h128C: out_word = 8'hDF;
		16'h128D: out_word = 8'h0E;
		16'h128E: out_word = 8'hFD;
		16'h128F: out_word = 8'h36;
		16'h1290: out_word = 8'h31;
		16'h1291: out_word = 8'h02;
		16'h1292: out_word = 8'hCD;
		16'h1293: out_word = 8'h6B;
		16'h1294: out_word = 8'h0D;
		16'h1295: out_word = 8'hAF;
		16'h1296: out_word = 8'h11;
		16'h1297: out_word = 8'h38;
		16'h1298: out_word = 8'h15;
		16'h1299: out_word = 8'hCD;
		16'h129A: out_word = 8'h0A;
		16'h129B: out_word = 8'h0C;
		16'h129C: out_word = 8'hFD;
		16'h129D: out_word = 8'hCB;
		16'h129E: out_word = 8'h02;
		16'h129F: out_word = 8'hEE;
		16'h12A0: out_word = 8'h18;
		16'h12A1: out_word = 8'h07;
		16'h12A2: out_word = 8'hFD;
		16'h12A3: out_word = 8'h36;
		16'h12A4: out_word = 8'h31;
		16'h12A5: out_word = 8'h02;
		16'h12A6: out_word = 8'hCD;
		16'h12A7: out_word = 8'h95;
		16'h12A8: out_word = 8'h17;
		16'h12A9: out_word = 8'hCD;
		16'h12AA: out_word = 8'hB0;
		16'h12AB: out_word = 8'h16;
		16'h12AC: out_word = 8'h3E;
		16'h12AD: out_word = 8'h00;
		16'h12AE: out_word = 8'hCD;
		16'h12AF: out_word = 8'h01;
		16'h12B0: out_word = 8'h16;
		16'h12B1: out_word = 8'hCD;
		16'h12B2: out_word = 8'h2C;
		16'h12B3: out_word = 8'h0F;
		16'h12B4: out_word = 8'hCD;
		16'h12B5: out_word = 8'h17;
		16'h12B6: out_word = 8'h1B;
		16'h12B7: out_word = 8'hFD;
		16'h12B8: out_word = 8'hCB;
		16'h12B9: out_word = 8'h00;
		16'h12BA: out_word = 8'h7E;
		16'h12BB: out_word = 8'h20;
		16'h12BC: out_word = 8'h12;
		16'h12BD: out_word = 8'hFD;
		16'h12BE: out_word = 8'hCB;
		16'h12BF: out_word = 8'h30;
		16'h12C0: out_word = 8'h66;
		16'h12C1: out_word = 8'h28;
		16'h12C2: out_word = 8'h40;
		16'h12C3: out_word = 8'h2A;
		16'h12C4: out_word = 8'h59;
		16'h12C5: out_word = 8'h5C;
		16'h12C6: out_word = 8'hCD;
		16'h12C7: out_word = 8'hA7;
		16'h12C8: out_word = 8'h11;
		16'h12C9: out_word = 8'hFD;
		16'h12CA: out_word = 8'h36;
		16'h12CB: out_word = 8'h00;
		16'h12CC: out_word = 8'hFF;
		16'h12CD: out_word = 8'h18;
		16'h12CE: out_word = 8'hDD;
		16'h12CF: out_word = 8'h2A;
		16'h12D0: out_word = 8'h59;
		16'h12D1: out_word = 8'h5C;
		16'h12D2: out_word = 8'h22;
		16'h12D3: out_word = 8'h5D;
		16'h12D4: out_word = 8'h5C;
		16'h12D5: out_word = 8'hCD;
		16'h12D6: out_word = 8'hFB;
		16'h12D7: out_word = 8'h19;
		16'h12D8: out_word = 8'h78;
		16'h12D9: out_word = 8'hB1;
		16'h12DA: out_word = 8'hC2;
		16'h12DB: out_word = 8'h5D;
		16'h12DC: out_word = 8'h15;
		16'h12DD: out_word = 8'hDF;
		16'h12DE: out_word = 8'hFE;
		16'h12DF: out_word = 8'h0D;
		16'h12E0: out_word = 8'h28;
		16'h12E1: out_word = 8'hC0;
		16'h12E2: out_word = 8'hFD;
		16'h12E3: out_word = 8'hCB;
		16'h12E4: out_word = 8'h30;
		16'h12E5: out_word = 8'h46;
		16'h12E6: out_word = 8'hC4;
		16'h12E7: out_word = 8'hAF;
		16'h12E8: out_word = 8'h0D;
		16'h12E9: out_word = 8'hCD;
		16'h12EA: out_word = 8'h6E;
		16'h12EB: out_word = 8'h0D;
		16'h12EC: out_word = 8'h3E;
		16'h12ED: out_word = 8'h19;
		16'h12EE: out_word = 8'hFD;
		16'h12EF: out_word = 8'h96;
		16'h12F0: out_word = 8'h4F;
		16'h12F1: out_word = 8'h32;
		16'h12F2: out_word = 8'h8C;
		16'h12F3: out_word = 8'h5C;
		16'h12F4: out_word = 8'hFD;
		16'h12F5: out_word = 8'hCB;
		16'h12F6: out_word = 8'h01;
		16'h12F7: out_word = 8'hFE;
		16'h12F8: out_word = 8'hFD;
		16'h12F9: out_word = 8'h36;
		16'h12FA: out_word = 8'h00;
		16'h12FB: out_word = 8'hFF;
		16'h12FC: out_word = 8'hFD;
		16'h12FD: out_word = 8'h36;
		16'h12FE: out_word = 8'h0A;
		16'h12FF: out_word = 8'h01;
		16'h1300: out_word = 8'hCD;
		16'h1301: out_word = 8'h8A;
		16'h1302: out_word = 8'h1B;
		16'h1303: out_word = 8'h76;
		16'h1304: out_word = 8'hFD;
		16'h1305: out_word = 8'hCB;
		16'h1306: out_word = 8'h01;
		16'h1307: out_word = 8'hAE;
		16'h1308: out_word = 8'hFD;
		16'h1309: out_word = 8'hCB;
		16'h130A: out_word = 8'h30;
		16'h130B: out_word = 8'h4E;
		16'h130C: out_word = 8'hC4;
		16'h130D: out_word = 8'hCD;
		16'h130E: out_word = 8'h0E;
		16'h130F: out_word = 8'h3A;
		16'h1310: out_word = 8'h3A;
		16'h1311: out_word = 8'h5C;
		16'h1312: out_word = 8'h3C;
		16'h1313: out_word = 8'hF5;
		16'h1314: out_word = 8'h21;
		16'h1315: out_word = 8'h00;
		16'h1316: out_word = 8'h00;
		16'h1317: out_word = 8'hFD;
		16'h1318: out_word = 8'h74;
		16'h1319: out_word = 8'h37;
		16'h131A: out_word = 8'hFD;
		16'h131B: out_word = 8'h74;
		16'h131C: out_word = 8'h26;
		16'h131D: out_word = 8'h22;
		16'h131E: out_word = 8'h0B;
		16'h131F: out_word = 8'h5C;
		16'h1320: out_word = 8'h21;
		16'h1321: out_word = 8'h01;
		16'h1322: out_word = 8'h00;
		16'h1323: out_word = 8'h22;
		16'h1324: out_word = 8'h16;
		16'h1325: out_word = 8'h5C;
		16'h1326: out_word = 8'hCD;
		16'h1327: out_word = 8'hB0;
		16'h1328: out_word = 8'h16;
		16'h1329: out_word = 8'hFD;
		16'h132A: out_word = 8'hCB;
		16'h132B: out_word = 8'h37;
		16'h132C: out_word = 8'hAE;
		16'h132D: out_word = 8'hCD;
		16'h132E: out_word = 8'h6E;
		16'h132F: out_word = 8'h0D;
		16'h1330: out_word = 8'hFD;
		16'h1331: out_word = 8'hCB;
		16'h1332: out_word = 8'h02;
		16'h1333: out_word = 8'hEE;
		16'h1334: out_word = 8'hF1;
		16'h1335: out_word = 8'h47;
		16'h1336: out_word = 8'hFE;
		16'h1337: out_word = 8'h0A;
		16'h1338: out_word = 8'h38;
		16'h1339: out_word = 8'h02;
		16'h133A: out_word = 8'hC6;
		16'h133B: out_word = 8'h07;
		16'h133C: out_word = 8'hCD;
		16'h133D: out_word = 8'hEF;
		16'h133E: out_word = 8'h15;
		16'h133F: out_word = 8'h3E;
		16'h1340: out_word = 8'h20;
		16'h1341: out_word = 8'hD7;
		16'h1342: out_word = 8'h78;
		16'h1343: out_word = 8'h11;
		16'h1344: out_word = 8'h91;
		16'h1345: out_word = 8'h13;
		16'h1346: out_word = 8'hCD;
		16'h1347: out_word = 8'h0A;
		16'h1348: out_word = 8'h0C;
		16'h1349: out_word = 8'hCD;
		16'h134A: out_word = 8'h3B;
		16'h134B: out_word = 8'h3B;
		16'h134C: out_word = 8'h00;
		16'h134D: out_word = 8'hCD;
		16'h134E: out_word = 8'h0A;
		16'h134F: out_word = 8'h0C;
		16'h1350: out_word = 8'hED;
		16'h1351: out_word = 8'h4B;
		16'h1352: out_word = 8'h45;
		16'h1353: out_word = 8'h5C;
		16'h1354: out_word = 8'hCD;
		16'h1355: out_word = 8'h1B;
		16'h1356: out_word = 8'h1A;
		16'h1357: out_word = 8'h3E;
		16'h1358: out_word = 8'h3A;
		16'h1359: out_word = 8'hD7;
		16'h135A: out_word = 8'hFD;
		16'h135B: out_word = 8'h4E;
		16'h135C: out_word = 8'h0D;
		16'h135D: out_word = 8'h06;
		16'h135E: out_word = 8'h00;
		16'h135F: out_word = 8'hCD;
		16'h1360: out_word = 8'h1B;
		16'h1361: out_word = 8'h1A;
		16'h1362: out_word = 8'hCD;
		16'h1363: out_word = 8'h97;
		16'h1364: out_word = 8'h10;
		16'h1365: out_word = 8'h3A;
		16'h1366: out_word = 8'h3A;
		16'h1367: out_word = 8'h5C;
		16'h1368: out_word = 8'h3C;
		16'h1369: out_word = 8'h28;
		16'h136A: out_word = 8'h1B;
		16'h136B: out_word = 8'hFE;
		16'h136C: out_word = 8'h09;
		16'h136D: out_word = 8'h28;
		16'h136E: out_word = 8'h04;
		16'h136F: out_word = 8'hFE;
		16'h1370: out_word = 8'h15;
		16'h1371: out_word = 8'h20;
		16'h1372: out_word = 8'h03;
		16'h1373: out_word = 8'hFD;
		16'h1374: out_word = 8'h34;
		16'h1375: out_word = 8'h0D;
		16'h1376: out_word = 8'h01;
		16'h1377: out_word = 8'h03;
		16'h1378: out_word = 8'h00;
		16'h1379: out_word = 8'h11;
		16'h137A: out_word = 8'h70;
		16'h137B: out_word = 8'h5C;
		16'h137C: out_word = 8'h21;
		16'h137D: out_word = 8'h44;
		16'h137E: out_word = 8'h5C;
		16'h137F: out_word = 8'hCB;
		16'h1380: out_word = 8'h7E;
		16'h1381: out_word = 8'h28;
		16'h1382: out_word = 8'h01;
		16'h1383: out_word = 8'h09;
		16'h1384: out_word = 8'hED;
		16'h1385: out_word = 8'hB8;
		16'h1386: out_word = 8'hFD;
		16'h1387: out_word = 8'h36;
		16'h1388: out_word = 8'h0A;
		16'h1389: out_word = 8'hFF;
		16'h138A: out_word = 8'hFD;
		16'h138B: out_word = 8'hCB;
		16'h138C: out_word = 8'h01;
		16'h138D: out_word = 8'h9E;
		16'h138E: out_word = 8'hC3;
		16'h138F: out_word = 8'hAC;
		16'h1390: out_word = 8'h12;
		16'h1391: out_word = 8'h80;
		16'h1392: out_word = 8'h4F;
		16'h1393: out_word = 8'hCB;
		16'h1394: out_word = 8'h4E;
		16'h1395: out_word = 8'h45;
		16'h1396: out_word = 8'h58;
		16'h1397: out_word = 8'h54;
		16'h1398: out_word = 8'h20;
		16'h1399: out_word = 8'h77;
		16'h139A: out_word = 8'h69;
		16'h139B: out_word = 8'h74;
		16'h139C: out_word = 8'h68;
		16'h139D: out_word = 8'h6F;
		16'h139E: out_word = 8'h75;
		16'h139F: out_word = 8'h74;
		16'h13A0: out_word = 8'h20;
		16'h13A1: out_word = 8'h46;
		16'h13A2: out_word = 8'h4F;
		16'h13A3: out_word = 8'hD2;
		16'h13A4: out_word = 8'h56;
		16'h13A5: out_word = 8'h61;
		16'h13A6: out_word = 8'h72;
		16'h13A7: out_word = 8'h69;
		16'h13A8: out_word = 8'h61;
		16'h13A9: out_word = 8'h62;
		16'h13AA: out_word = 8'h6C;
		16'h13AB: out_word = 8'h65;
		16'h13AC: out_word = 8'h20;
		16'h13AD: out_word = 8'h6E;
		16'h13AE: out_word = 8'h6F;
		16'h13AF: out_word = 8'h74;
		16'h13B0: out_word = 8'h20;
		16'h13B1: out_word = 8'h66;
		16'h13B2: out_word = 8'h6F;
		16'h13B3: out_word = 8'h75;
		16'h13B4: out_word = 8'h6E;
		16'h13B5: out_word = 8'hE4;
		16'h13B6: out_word = 8'h53;
		16'h13B7: out_word = 8'h75;
		16'h13B8: out_word = 8'h62;
		16'h13B9: out_word = 8'h73;
		16'h13BA: out_word = 8'h63;
		16'h13BB: out_word = 8'h72;
		16'h13BC: out_word = 8'h69;
		16'h13BD: out_word = 8'h70;
		16'h13BE: out_word = 8'h74;
		16'h13BF: out_word = 8'h20;
		16'h13C0: out_word = 8'h77;
		16'h13C1: out_word = 8'h72;
		16'h13C2: out_word = 8'h6F;
		16'h13C3: out_word = 8'h6E;
		16'h13C4: out_word = 8'hE7;
		16'h13C5: out_word = 8'h4F;
		16'h13C6: out_word = 8'h75;
		16'h13C7: out_word = 8'h74;
		16'h13C8: out_word = 8'h20;
		16'h13C9: out_word = 8'h6F;
		16'h13CA: out_word = 8'h66;
		16'h13CB: out_word = 8'h20;
		16'h13CC: out_word = 8'h6D;
		16'h13CD: out_word = 8'h65;
		16'h13CE: out_word = 8'h6D;
		16'h13CF: out_word = 8'h6F;
		16'h13D0: out_word = 8'h72;
		16'h13D1: out_word = 8'hF9;
		16'h13D2: out_word = 8'h4F;
		16'h13D3: out_word = 8'h75;
		16'h13D4: out_word = 8'h74;
		16'h13D5: out_word = 8'h20;
		16'h13D6: out_word = 8'h6F;
		16'h13D7: out_word = 8'h66;
		16'h13D8: out_word = 8'h20;
		16'h13D9: out_word = 8'h73;
		16'h13DA: out_word = 8'h63;
		16'h13DB: out_word = 8'h72;
		16'h13DC: out_word = 8'h65;
		16'h13DD: out_word = 8'h65;
		16'h13DE: out_word = 8'hEE;
		16'h13DF: out_word = 8'h4E;
		16'h13E0: out_word = 8'h75;
		16'h13E1: out_word = 8'h6D;
		16'h13E2: out_word = 8'h62;
		16'h13E3: out_word = 8'h65;
		16'h13E4: out_word = 8'h72;
		16'h13E5: out_word = 8'h20;
		16'h13E6: out_word = 8'h74;
		16'h13E7: out_word = 8'h6F;
		16'h13E8: out_word = 8'h6F;
		16'h13E9: out_word = 8'h20;
		16'h13EA: out_word = 8'h62;
		16'h13EB: out_word = 8'h69;
		16'h13EC: out_word = 8'hE7;
		16'h13ED: out_word = 8'h52;
		16'h13EE: out_word = 8'h45;
		16'h13EF: out_word = 8'h54;
		16'h13F0: out_word = 8'h55;
		16'h13F1: out_word = 8'h52;
		16'h13F2: out_word = 8'h4E;
		16'h13F3: out_word = 8'h20;
		16'h13F4: out_word = 8'h77;
		16'h13F5: out_word = 8'h69;
		16'h13F6: out_word = 8'h74;
		16'h13F7: out_word = 8'h68;
		16'h13F8: out_word = 8'h6F;
		16'h13F9: out_word = 8'h75;
		16'h13FA: out_word = 8'h74;
		16'h13FB: out_word = 8'h20;
		16'h13FC: out_word = 8'h47;
		16'h13FD: out_word = 8'h4F;
		16'h13FE: out_word = 8'h53;
		16'h13FF: out_word = 8'h55;
		16'h1400: out_word = 8'hC2;
		16'h1401: out_word = 8'h45;
		16'h1402: out_word = 8'h6E;
		16'h1403: out_word = 8'h64;
		16'h1404: out_word = 8'h20;
		16'h1405: out_word = 8'h6F;
		16'h1406: out_word = 8'h66;
		16'h1407: out_word = 8'h20;
		16'h1408: out_word = 8'h66;
		16'h1409: out_word = 8'h69;
		16'h140A: out_word = 8'h6C;
		16'h140B: out_word = 8'hE5;
		16'h140C: out_word = 8'h53;
		16'h140D: out_word = 8'h54;
		16'h140E: out_word = 8'h4F;
		16'h140F: out_word = 8'h50;
		16'h1410: out_word = 8'h20;
		16'h1411: out_word = 8'h73;
		16'h1412: out_word = 8'h74;
		16'h1413: out_word = 8'h61;
		16'h1414: out_word = 8'h74;
		16'h1415: out_word = 8'h65;
		16'h1416: out_word = 8'h6D;
		16'h1417: out_word = 8'h65;
		16'h1418: out_word = 8'h6E;
		16'h1419: out_word = 8'hF4;
		16'h141A: out_word = 8'h49;
		16'h141B: out_word = 8'h6E;
		16'h141C: out_word = 8'h76;
		16'h141D: out_word = 8'h61;
		16'h141E: out_word = 8'h6C;
		16'h141F: out_word = 8'h69;
		16'h1420: out_word = 8'h64;
		16'h1421: out_word = 8'h20;
		16'h1422: out_word = 8'h61;
		16'h1423: out_word = 8'h72;
		16'h1424: out_word = 8'h67;
		16'h1425: out_word = 8'h75;
		16'h1426: out_word = 8'h6D;
		16'h1427: out_word = 8'h65;
		16'h1428: out_word = 8'h6E;
		16'h1429: out_word = 8'hF4;
		16'h142A: out_word = 8'h49;
		16'h142B: out_word = 8'h6E;
		16'h142C: out_word = 8'h74;
		16'h142D: out_word = 8'h65;
		16'h142E: out_word = 8'h67;
		16'h142F: out_word = 8'h65;
		16'h1430: out_word = 8'h72;
		16'h1431: out_word = 8'h20;
		16'h1432: out_word = 8'h6F;
		16'h1433: out_word = 8'h75;
		16'h1434: out_word = 8'h74;
		16'h1435: out_word = 8'h20;
		16'h1436: out_word = 8'h6F;
		16'h1437: out_word = 8'h66;
		16'h1438: out_word = 8'h20;
		16'h1439: out_word = 8'h72;
		16'h143A: out_word = 8'h61;
		16'h143B: out_word = 8'h6E;
		16'h143C: out_word = 8'h67;
		16'h143D: out_word = 8'hE5;
		16'h143E: out_word = 8'h4E;
		16'h143F: out_word = 8'h6F;
		16'h1440: out_word = 8'h6E;
		16'h1441: out_word = 8'h73;
		16'h1442: out_word = 8'h65;
		16'h1443: out_word = 8'h6E;
		16'h1444: out_word = 8'h73;
		16'h1445: out_word = 8'h65;
		16'h1446: out_word = 8'h20;
		16'h1447: out_word = 8'h69;
		16'h1448: out_word = 8'h6E;
		16'h1449: out_word = 8'h20;
		16'h144A: out_word = 8'h42;
		16'h144B: out_word = 8'h41;
		16'h144C: out_word = 8'h53;
		16'h144D: out_word = 8'h49;
		16'h144E: out_word = 8'hC3;
		16'h144F: out_word = 8'h42;
		16'h1450: out_word = 8'h52;
		16'h1451: out_word = 8'h45;
		16'h1452: out_word = 8'h41;
		16'h1453: out_word = 8'h4B;
		16'h1454: out_word = 8'h20;
		16'h1455: out_word = 8'h2D;
		16'h1456: out_word = 8'h20;
		16'h1457: out_word = 8'h43;
		16'h1458: out_word = 8'h4F;
		16'h1459: out_word = 8'h4E;
		16'h145A: out_word = 8'h54;
		16'h145B: out_word = 8'h20;
		16'h145C: out_word = 8'h72;
		16'h145D: out_word = 8'h65;
		16'h145E: out_word = 8'h70;
		16'h145F: out_word = 8'h65;
		16'h1460: out_word = 8'h61;
		16'h1461: out_word = 8'h74;
		16'h1462: out_word = 8'hF3;
		16'h1463: out_word = 8'h4F;
		16'h1464: out_word = 8'h75;
		16'h1465: out_word = 8'h74;
		16'h1466: out_word = 8'h20;
		16'h1467: out_word = 8'h6F;
		16'h1468: out_word = 8'h66;
		16'h1469: out_word = 8'h20;
		16'h146A: out_word = 8'h44;
		16'h146B: out_word = 8'h41;
		16'h146C: out_word = 8'h54;
		16'h146D: out_word = 8'hC1;
		16'h146E: out_word = 8'h49;
		16'h146F: out_word = 8'h6E;
		16'h1470: out_word = 8'h76;
		16'h1471: out_word = 8'h61;
		16'h1472: out_word = 8'h6C;
		16'h1473: out_word = 8'h69;
		16'h1474: out_word = 8'h64;
		16'h1475: out_word = 8'h20;
		16'h1476: out_word = 8'h66;
		16'h1477: out_word = 8'h69;
		16'h1478: out_word = 8'h6C;
		16'h1479: out_word = 8'h65;
		16'h147A: out_word = 8'h20;
		16'h147B: out_word = 8'h6E;
		16'h147C: out_word = 8'h61;
		16'h147D: out_word = 8'h6D;
		16'h147E: out_word = 8'hE5;
		16'h147F: out_word = 8'h4E;
		16'h1480: out_word = 8'h6F;
		16'h1481: out_word = 8'h20;
		16'h1482: out_word = 8'h72;
		16'h1483: out_word = 8'h6F;
		16'h1484: out_word = 8'h6F;
		16'h1485: out_word = 8'h6D;
		16'h1486: out_word = 8'h20;
		16'h1487: out_word = 8'h66;
		16'h1488: out_word = 8'h6F;
		16'h1489: out_word = 8'h72;
		16'h148A: out_word = 8'h20;
		16'h148B: out_word = 8'h6C;
		16'h148C: out_word = 8'h69;
		16'h148D: out_word = 8'h6E;
		16'h148E: out_word = 8'hE5;
		16'h148F: out_word = 8'h53;
		16'h1490: out_word = 8'h54;
		16'h1491: out_word = 8'h4F;
		16'h1492: out_word = 8'h50;
		16'h1493: out_word = 8'h20;
		16'h1494: out_word = 8'h69;
		16'h1495: out_word = 8'h6E;
		16'h1496: out_word = 8'h20;
		16'h1497: out_word = 8'h49;
		16'h1498: out_word = 8'h4E;
		16'h1499: out_word = 8'h50;
		16'h149A: out_word = 8'h55;
		16'h149B: out_word = 8'hD4;
		16'h149C: out_word = 8'h46;
		16'h149D: out_word = 8'h4F;
		16'h149E: out_word = 8'h52;
		16'h149F: out_word = 8'h20;
		16'h14A0: out_word = 8'h77;
		16'h14A1: out_word = 8'h69;
		16'h14A2: out_word = 8'h74;
		16'h14A3: out_word = 8'h68;
		16'h14A4: out_word = 8'h6F;
		16'h14A5: out_word = 8'h75;
		16'h14A6: out_word = 8'h74;
		16'h14A7: out_word = 8'h20;
		16'h14A8: out_word = 8'h4E;
		16'h14A9: out_word = 8'h45;
		16'h14AA: out_word = 8'h58;
		16'h14AB: out_word = 8'hD4;
		16'h14AC: out_word = 8'h49;
		16'h14AD: out_word = 8'h6E;
		16'h14AE: out_word = 8'h76;
		16'h14AF: out_word = 8'h61;
		16'h14B0: out_word = 8'h6C;
		16'h14B1: out_word = 8'h69;
		16'h14B2: out_word = 8'h64;
		16'h14B3: out_word = 8'h20;
		16'h14B4: out_word = 8'h49;
		16'h14B5: out_word = 8'h2F;
		16'h14B6: out_word = 8'h4F;
		16'h14B7: out_word = 8'h20;
		16'h14B8: out_word = 8'h64;
		16'h14B9: out_word = 8'h65;
		16'h14BA: out_word = 8'h76;
		16'h14BB: out_word = 8'h69;
		16'h14BC: out_word = 8'h63;
		16'h14BD: out_word = 8'hE5;
		16'h14BE: out_word = 8'h49;
		16'h14BF: out_word = 8'h6E;
		16'h14C0: out_word = 8'h76;
		16'h14C1: out_word = 8'h61;
		16'h14C2: out_word = 8'h6C;
		16'h14C3: out_word = 8'h69;
		16'h14C4: out_word = 8'h64;
		16'h14C5: out_word = 8'h20;
		16'h14C6: out_word = 8'h63;
		16'h14C7: out_word = 8'h6F;
		16'h14C8: out_word = 8'h6C;
		16'h14C9: out_word = 8'h6F;
		16'h14CA: out_word = 8'h75;
		16'h14CB: out_word = 8'hF2;
		16'h14CC: out_word = 8'h42;
		16'h14CD: out_word = 8'h52;
		16'h14CE: out_word = 8'h45;
		16'h14CF: out_word = 8'h41;
		16'h14D0: out_word = 8'h4B;
		16'h14D1: out_word = 8'h20;
		16'h14D2: out_word = 8'h69;
		16'h14D3: out_word = 8'h6E;
		16'h14D4: out_word = 8'h74;
		16'h14D5: out_word = 8'h6F;
		16'h14D6: out_word = 8'h20;
		16'h14D7: out_word = 8'h70;
		16'h14D8: out_word = 8'h72;
		16'h14D9: out_word = 8'h6F;
		16'h14DA: out_word = 8'h67;
		16'h14DB: out_word = 8'h72;
		16'h14DC: out_word = 8'h61;
		16'h14DD: out_word = 8'hED;
		16'h14DE: out_word = 8'h52;
		16'h14DF: out_word = 8'h41;
		16'h14E0: out_word = 8'h4D;
		16'h14E1: out_word = 8'h54;
		16'h14E2: out_word = 8'h4F;
		16'h14E3: out_word = 8'h50;
		16'h14E4: out_word = 8'h20;
		16'h14E5: out_word = 8'h6E;
		16'h14E6: out_word = 8'h6F;
		16'h14E7: out_word = 8'h20;
		16'h14E8: out_word = 8'h67;
		16'h14E9: out_word = 8'h6F;
		16'h14EA: out_word = 8'h6F;
		16'h14EB: out_word = 8'hE4;
		16'h14EC: out_word = 8'h53;
		16'h14ED: out_word = 8'h74;
		16'h14EE: out_word = 8'h61;
		16'h14EF: out_word = 8'h74;
		16'h14F0: out_word = 8'h65;
		16'h14F1: out_word = 8'h6D;
		16'h14F2: out_word = 8'h65;
		16'h14F3: out_word = 8'h6E;
		16'h14F4: out_word = 8'h74;
		16'h14F5: out_word = 8'h20;
		16'h14F6: out_word = 8'h6C;
		16'h14F7: out_word = 8'h6F;
		16'h14F8: out_word = 8'h73;
		16'h14F9: out_word = 8'hF4;
		16'h14FA: out_word = 8'h49;
		16'h14FB: out_word = 8'h6E;
		16'h14FC: out_word = 8'h76;
		16'h14FD: out_word = 8'h61;
		16'h14FE: out_word = 8'h6C;
		16'h14FF: out_word = 8'h69;
		16'h1500: out_word = 8'h64;
		16'h1501: out_word = 8'h20;
		16'h1502: out_word = 8'h73;
		16'h1503: out_word = 8'h74;
		16'h1504: out_word = 8'h72;
		16'h1505: out_word = 8'h65;
		16'h1506: out_word = 8'h61;
		16'h1507: out_word = 8'hED;
		16'h1508: out_word = 8'h46;
		16'h1509: out_word = 8'h4E;
		16'h150A: out_word = 8'h20;
		16'h150B: out_word = 8'h77;
		16'h150C: out_word = 8'h69;
		16'h150D: out_word = 8'h74;
		16'h150E: out_word = 8'h68;
		16'h150F: out_word = 8'h6F;
		16'h1510: out_word = 8'h75;
		16'h1511: out_word = 8'h74;
		16'h1512: out_word = 8'h20;
		16'h1513: out_word = 8'h44;
		16'h1514: out_word = 8'h45;
		16'h1515: out_word = 8'hC6;
		16'h1516: out_word = 8'h50;
		16'h1517: out_word = 8'h61;
		16'h1518: out_word = 8'h72;
		16'h1519: out_word = 8'h61;
		16'h151A: out_word = 8'h6D;
		16'h151B: out_word = 8'h65;
		16'h151C: out_word = 8'h74;
		16'h151D: out_word = 8'h65;
		16'h151E: out_word = 8'h72;
		16'h151F: out_word = 8'h20;
		16'h1520: out_word = 8'h65;
		16'h1521: out_word = 8'h72;
		16'h1522: out_word = 8'h72;
		16'h1523: out_word = 8'h6F;
		16'h1524: out_word = 8'hF2;
		16'h1525: out_word = 8'h54;
		16'h1526: out_word = 8'h61;
		16'h1527: out_word = 8'h70;
		16'h1528: out_word = 8'h65;
		16'h1529: out_word = 8'h20;
		16'h152A: out_word = 8'h6C;
		16'h152B: out_word = 8'h6F;
		16'h152C: out_word = 8'h61;
		16'h152D: out_word = 8'h64;
		16'h152E: out_word = 8'h69;
		16'h152F: out_word = 8'h6E;
		16'h1530: out_word = 8'h67;
		16'h1531: out_word = 8'h20;
		16'h1532: out_word = 8'h65;
		16'h1533: out_word = 8'h72;
		16'h1534: out_word = 8'h72;
		16'h1535: out_word = 8'h6F;
		16'h1536: out_word = 8'hF2;
		16'h1537: out_word = 8'h2C;
		16'h1538: out_word = 8'hA0;
		16'h1539: out_word = 8'h7F;
		16'h153A: out_word = 8'h20;
		16'h153B: out_word = 8'h31;
		16'h153C: out_word = 8'h39;
		16'h153D: out_word = 8'h38;
		16'h153E: out_word = 8'h32;
		16'h153F: out_word = 8'h20;
		16'h1540: out_word = 8'h53;
		16'h1541: out_word = 8'h69;
		16'h1542: out_word = 8'h6E;
		16'h1543: out_word = 8'h63;
		16'h1544: out_word = 8'h6C;
		16'h1545: out_word = 8'h61;
		16'h1546: out_word = 8'h69;
		16'h1547: out_word = 8'h72;
		16'h1548: out_word = 8'h20;
		16'h1549: out_word = 8'h52;
		16'h154A: out_word = 8'h65;
		16'h154B: out_word = 8'h73;
		16'h154C: out_word = 8'h65;
		16'h154D: out_word = 8'h61;
		16'h154E: out_word = 8'h72;
		16'h154F: out_word = 8'h63;
		16'h1550: out_word = 8'h68;
		16'h1551: out_word = 8'h20;
		16'h1552: out_word = 8'h4C;
		16'h1553: out_word = 8'h74;
		16'h1554: out_word = 8'hE4;
		16'h1555: out_word = 8'h3E;
		16'h1556: out_word = 8'h10;
		16'h1557: out_word = 8'h01;
		16'h1558: out_word = 8'h00;
		16'h1559: out_word = 8'h00;
		16'h155A: out_word = 8'hC3;
		16'h155B: out_word = 8'h13;
		16'h155C: out_word = 8'h13;
		16'h155D: out_word = 8'hED;
		16'h155E: out_word = 8'h43;
		16'h155F: out_word = 8'h49;
		16'h1560: out_word = 8'h5C;
		16'h1561: out_word = 8'h2A;
		16'h1562: out_word = 8'h5D;
		16'h1563: out_word = 8'h5C;
		16'h1564: out_word = 8'hEB;
		16'h1565: out_word = 8'h21;
		16'h1566: out_word = 8'h55;
		16'h1567: out_word = 8'h15;
		16'h1568: out_word = 8'hE5;
		16'h1569: out_word = 8'h2A;
		16'h156A: out_word = 8'h61;
		16'h156B: out_word = 8'h5C;
		16'h156C: out_word = 8'h37;
		16'h156D: out_word = 8'hED;
		16'h156E: out_word = 8'h52;
		16'h156F: out_word = 8'hE5;
		16'h1570: out_word = 8'h60;
		16'h1571: out_word = 8'h69;
		16'h1572: out_word = 8'hCD;
		16'h1573: out_word = 8'h6E;
		16'h1574: out_word = 8'h19;
		16'h1575: out_word = 8'h20;
		16'h1576: out_word = 8'h06;
		16'h1577: out_word = 8'hCD;
		16'h1578: out_word = 8'hB8;
		16'h1579: out_word = 8'h19;
		16'h157A: out_word = 8'hCD;
		16'h157B: out_word = 8'hE8;
		16'h157C: out_word = 8'h19;
		16'h157D: out_word = 8'hC1;
		16'h157E: out_word = 8'h79;
		16'h157F: out_word = 8'h3D;
		16'h1580: out_word = 8'hB0;
		16'h1581: out_word = 8'h28;
		16'h1582: out_word = 8'h28;
		16'h1583: out_word = 8'hC5;
		16'h1584: out_word = 8'h03;
		16'h1585: out_word = 8'h03;
		16'h1586: out_word = 8'h03;
		16'h1587: out_word = 8'h03;
		16'h1588: out_word = 8'h2B;
		16'h1589: out_word = 8'hED;
		16'h158A: out_word = 8'h5B;
		16'h158B: out_word = 8'h53;
		16'h158C: out_word = 8'h5C;
		16'h158D: out_word = 8'hD5;
		16'h158E: out_word = 8'hCD;
		16'h158F: out_word = 8'h55;
		16'h1590: out_word = 8'h16;
		16'h1591: out_word = 8'hE1;
		16'h1592: out_word = 8'h22;
		16'h1593: out_word = 8'h53;
		16'h1594: out_word = 8'h5C;
		16'h1595: out_word = 8'hC1;
		16'h1596: out_word = 8'hC5;
		16'h1597: out_word = 8'h13;
		16'h1598: out_word = 8'h2A;
		16'h1599: out_word = 8'h61;
		16'h159A: out_word = 8'h5C;
		16'h159B: out_word = 8'h2B;
		16'h159C: out_word = 8'h2B;
		16'h159D: out_word = 8'hED;
		16'h159E: out_word = 8'hB8;
		16'h159F: out_word = 8'h2A;
		16'h15A0: out_word = 8'h49;
		16'h15A1: out_word = 8'h5C;
		16'h15A2: out_word = 8'hEB;
		16'h15A3: out_word = 8'hC1;
		16'h15A4: out_word = 8'h70;
		16'h15A5: out_word = 8'h2B;
		16'h15A6: out_word = 8'h71;
		16'h15A7: out_word = 8'h2B;
		16'h15A8: out_word = 8'h73;
		16'h15A9: out_word = 8'h2B;
		16'h15AA: out_word = 8'h72;
		16'h15AB: out_word = 8'hF1;
		16'h15AC: out_word = 8'hC3;
		16'h15AD: out_word = 8'hA2;
		16'h15AE: out_word = 8'h12;
		16'h15AF: out_word = 8'hF4;
		16'h15B0: out_word = 8'h09;
		16'h15B1: out_word = 8'hA8;
		16'h15B2: out_word = 8'h10;
		16'h15B3: out_word = 8'h4B;
		16'h15B4: out_word = 8'hF4;
		16'h15B5: out_word = 8'h09;
		16'h15B6: out_word = 8'hC4;
		16'h15B7: out_word = 8'h15;
		16'h15B8: out_word = 8'h53;
		16'h15B9: out_word = 8'h81;
		16'h15BA: out_word = 8'h0F;
		16'h15BB: out_word = 8'hC4;
		16'h15BC: out_word = 8'h15;
		16'h15BD: out_word = 8'h52;
		16'h15BE: out_word = 8'hF4;
		16'h15BF: out_word = 8'h09;
		16'h15C0: out_word = 8'hC4;
		16'h15C1: out_word = 8'h15;
		16'h15C2: out_word = 8'h50;
		16'h15C3: out_word = 8'h80;
		16'h15C4: out_word = 8'hCF;
		16'h15C5: out_word = 8'h12;
		16'h15C6: out_word = 8'h01;
		16'h15C7: out_word = 8'h00;
		16'h15C8: out_word = 8'h06;
		16'h15C9: out_word = 8'h00;
		16'h15CA: out_word = 8'h0B;
		16'h15CB: out_word = 8'h00;
		16'h15CC: out_word = 8'h01;
		16'h15CD: out_word = 8'h00;
		16'h15CE: out_word = 8'h01;
		16'h15CF: out_word = 8'h00;
		16'h15D0: out_word = 8'h06;
		16'h15D1: out_word = 8'h00;
		16'h15D2: out_word = 8'h10;
		16'h15D3: out_word = 8'h00;
		16'h15D4: out_word = 8'hFD;
		16'h15D5: out_word = 8'hCB;
		16'h15D6: out_word = 8'h02;
		16'h15D7: out_word = 8'h6E;
		16'h15D8: out_word = 8'h20;
		16'h15D9: out_word = 8'h04;
		16'h15DA: out_word = 8'hFD;
		16'h15DB: out_word = 8'hCB;
		16'h15DC: out_word = 8'h02;
		16'h15DD: out_word = 8'hDE;
		16'h15DE: out_word = 8'hCD;
		16'h15DF: out_word = 8'hE6;
		16'h15E0: out_word = 8'h15;
		16'h15E1: out_word = 8'hD8;
		16'h15E2: out_word = 8'h28;
		16'h15E3: out_word = 8'hFA;
		16'h15E4: out_word = 8'hCF;
		16'h15E5: out_word = 8'h07;
		16'h15E6: out_word = 8'hD9;
		16'h15E7: out_word = 8'hE5;
		16'h15E8: out_word = 8'h2A;
		16'h15E9: out_word = 8'h51;
		16'h15EA: out_word = 8'h5C;
		16'h15EB: out_word = 8'h23;
		16'h15EC: out_word = 8'h23;
		16'h15ED: out_word = 8'h18;
		16'h15EE: out_word = 8'h08;
		16'h15EF: out_word = 8'h1E;
		16'h15F0: out_word = 8'h30;
		16'h15F1: out_word = 8'h83;
		16'h15F2: out_word = 8'hD9;
		16'h15F3: out_word = 8'hE5;
		16'h15F4: out_word = 8'h2A;
		16'h15F5: out_word = 8'h51;
		16'h15F6: out_word = 8'h5C;
		16'h15F7: out_word = 8'h5E;
		16'h15F8: out_word = 8'h23;
		16'h15F9: out_word = 8'h56;
		16'h15FA: out_word = 8'hEB;
		16'h15FB: out_word = 8'hCD;
		16'h15FC: out_word = 8'h2C;
		16'h15FD: out_word = 8'h16;
		16'h15FE: out_word = 8'hE1;
		16'h15FF: out_word = 8'hD9;
		16'h1600: out_word = 8'hC9;
		16'h1601: out_word = 8'h87;
		16'h1602: out_word = 8'hC6;
		16'h1603: out_word = 8'h16;
		16'h1604: out_word = 8'h6F;
		16'h1605: out_word = 8'h26;
		16'h1606: out_word = 8'h5C;
		16'h1607: out_word = 8'h5E;
		16'h1608: out_word = 8'h23;
		16'h1609: out_word = 8'h56;
		16'h160A: out_word = 8'h7A;
		16'h160B: out_word = 8'hB3;
		16'h160C: out_word = 8'h20;
		16'h160D: out_word = 8'h02;
		16'h160E: out_word = 8'hCF;
		16'h160F: out_word = 8'h17;
		16'h1610: out_word = 8'h1B;
		16'h1611: out_word = 8'h2A;
		16'h1612: out_word = 8'h4F;
		16'h1613: out_word = 8'h5C;
		16'h1614: out_word = 8'h19;
		16'h1615: out_word = 8'h22;
		16'h1616: out_word = 8'h51;
		16'h1617: out_word = 8'h5C;
		16'h1618: out_word = 8'hFD;
		16'h1619: out_word = 8'hCB;
		16'h161A: out_word = 8'h30;
		16'h161B: out_word = 8'hA6;
		16'h161C: out_word = 8'h23;
		16'h161D: out_word = 8'h23;
		16'h161E: out_word = 8'h23;
		16'h161F: out_word = 8'h23;
		16'h1620: out_word = 8'h4E;
		16'h1621: out_word = 8'h21;
		16'h1622: out_word = 8'h2D;
		16'h1623: out_word = 8'h16;
		16'h1624: out_word = 8'hCD;
		16'h1625: out_word = 8'hDC;
		16'h1626: out_word = 8'h16;
		16'h1627: out_word = 8'hD0;
		16'h1628: out_word = 8'h16;
		16'h1629: out_word = 8'h00;
		16'h162A: out_word = 8'h5E;
		16'h162B: out_word = 8'h19;
		16'h162C: out_word = 8'hE9;
		16'h162D: out_word = 8'h4B;
		16'h162E: out_word = 8'h06;
		16'h162F: out_word = 8'h53;
		16'h1630: out_word = 8'h12;
		16'h1631: out_word = 8'h50;
		16'h1632: out_word = 8'h1B;
		16'h1633: out_word = 8'h00;
		16'h1634: out_word = 8'hFD;
		16'h1635: out_word = 8'hCB;
		16'h1636: out_word = 8'h02;
		16'h1637: out_word = 8'hC6;
		16'h1638: out_word = 8'hFD;
		16'h1639: out_word = 8'hCB;
		16'h163A: out_word = 8'h01;
		16'h163B: out_word = 8'hAE;
		16'h163C: out_word = 8'hFD;
		16'h163D: out_word = 8'hCB;
		16'h163E: out_word = 8'h30;
		16'h163F: out_word = 8'hE6;
		16'h1640: out_word = 8'h18;
		16'h1641: out_word = 8'h04;
		16'h1642: out_word = 8'hFD;
		16'h1643: out_word = 8'hCB;
		16'h1644: out_word = 8'h02;
		16'h1645: out_word = 8'h86;
		16'h1646: out_word = 8'hFD;
		16'h1647: out_word = 8'hCB;
		16'h1648: out_word = 8'h01;
		16'h1649: out_word = 8'h8E;
		16'h164A: out_word = 8'hC3;
		16'h164B: out_word = 8'h4D;
		16'h164C: out_word = 8'h0D;
		16'h164D: out_word = 8'hFD;
		16'h164E: out_word = 8'hCB;
		16'h164F: out_word = 8'h01;
		16'h1650: out_word = 8'hCE;
		16'h1651: out_word = 8'hC9;
		16'h1652: out_word = 8'h01;
		16'h1653: out_word = 8'h01;
		16'h1654: out_word = 8'h00;
		16'h1655: out_word = 8'hE5;
		16'h1656: out_word = 8'hCD;
		16'h1657: out_word = 8'h05;
		16'h1658: out_word = 8'h1F;
		16'h1659: out_word = 8'hE1;
		16'h165A: out_word = 8'hCD;
		16'h165B: out_word = 8'h64;
		16'h165C: out_word = 8'h16;
		16'h165D: out_word = 8'h2A;
		16'h165E: out_word = 8'h65;
		16'h165F: out_word = 8'h5C;
		16'h1660: out_word = 8'hEB;
		16'h1661: out_word = 8'hED;
		16'h1662: out_word = 8'hB8;
		16'h1663: out_word = 8'hC9;
		16'h1664: out_word = 8'hF5;
		16'h1665: out_word = 8'hE5;
		16'h1666: out_word = 8'h21;
		16'h1667: out_word = 8'h4B;
		16'h1668: out_word = 8'h5C;
		16'h1669: out_word = 8'h3E;
		16'h166A: out_word = 8'h0E;
		16'h166B: out_word = 8'h5E;
		16'h166C: out_word = 8'h23;
		16'h166D: out_word = 8'h56;
		16'h166E: out_word = 8'hE3;
		16'h166F: out_word = 8'hA7;
		16'h1670: out_word = 8'hED;
		16'h1671: out_word = 8'h52;
		16'h1672: out_word = 8'h19;
		16'h1673: out_word = 8'hE3;
		16'h1674: out_word = 8'h30;
		16'h1675: out_word = 8'h09;
		16'h1676: out_word = 8'hD5;
		16'h1677: out_word = 8'hEB;
		16'h1678: out_word = 8'h09;
		16'h1679: out_word = 8'hEB;
		16'h167A: out_word = 8'h72;
		16'h167B: out_word = 8'h2B;
		16'h167C: out_word = 8'h73;
		16'h167D: out_word = 8'h23;
		16'h167E: out_word = 8'hD1;
		16'h167F: out_word = 8'h23;
		16'h1680: out_word = 8'h3D;
		16'h1681: out_word = 8'h20;
		16'h1682: out_word = 8'hE8;
		16'h1683: out_word = 8'hEB;
		16'h1684: out_word = 8'hD1;
		16'h1685: out_word = 8'hF1;
		16'h1686: out_word = 8'hA7;
		16'h1687: out_word = 8'hED;
		16'h1688: out_word = 8'h52;
		16'h1689: out_word = 8'h44;
		16'h168A: out_word = 8'h4D;
		16'h168B: out_word = 8'h03;
		16'h168C: out_word = 8'h19;
		16'h168D: out_word = 8'hEB;
		16'h168E: out_word = 8'hC9;
		16'h168F: out_word = 8'h00;
		16'h1690: out_word = 8'h00;
		16'h1691: out_word = 8'hEB;
		16'h1692: out_word = 8'h11;
		16'h1693: out_word = 8'h8F;
		16'h1694: out_word = 8'h16;
		16'h1695: out_word = 8'h7E;
		16'h1696: out_word = 8'hE6;
		16'h1697: out_word = 8'hC0;
		16'h1698: out_word = 8'h20;
		16'h1699: out_word = 8'hF7;
		16'h169A: out_word = 8'h56;
		16'h169B: out_word = 8'h23;
		16'h169C: out_word = 8'h5E;
		16'h169D: out_word = 8'hC9;
		16'h169E: out_word = 8'h2A;
		16'h169F: out_word = 8'h63;
		16'h16A0: out_word = 8'h5C;
		16'h16A1: out_word = 8'h2B;
		16'h16A2: out_word = 8'hCD;
		16'h16A3: out_word = 8'h55;
		16'h16A4: out_word = 8'h16;
		16'h16A5: out_word = 8'h23;
		16'h16A6: out_word = 8'h23;
		16'h16A7: out_word = 8'hC1;
		16'h16A8: out_word = 8'hED;
		16'h16A9: out_word = 8'h43;
		16'h16AA: out_word = 8'h61;
		16'h16AB: out_word = 8'h5C;
		16'h16AC: out_word = 8'hC1;
		16'h16AD: out_word = 8'hEB;
		16'h16AE: out_word = 8'h23;
		16'h16AF: out_word = 8'hC9;
		16'h16B0: out_word = 8'h2A;
		16'h16B1: out_word = 8'h59;
		16'h16B2: out_word = 8'h5C;
		16'h16B3: out_word = 8'h36;
		16'h16B4: out_word = 8'h0D;
		16'h16B5: out_word = 8'h22;
		16'h16B6: out_word = 8'h5B;
		16'h16B7: out_word = 8'h5C;
		16'h16B8: out_word = 8'h23;
		16'h16B9: out_word = 8'h36;
		16'h16BA: out_word = 8'h80;
		16'h16BB: out_word = 8'h23;
		16'h16BC: out_word = 8'h22;
		16'h16BD: out_word = 8'h61;
		16'h16BE: out_word = 8'h5C;
		16'h16BF: out_word = 8'h2A;
		16'h16C0: out_word = 8'h61;
		16'h16C1: out_word = 8'h5C;
		16'h16C2: out_word = 8'h22;
		16'h16C3: out_word = 8'h63;
		16'h16C4: out_word = 8'h5C;
		16'h16C5: out_word = 8'h2A;
		16'h16C6: out_word = 8'h63;
		16'h16C7: out_word = 8'h5C;
		16'h16C8: out_word = 8'h22;
		16'h16C9: out_word = 8'h65;
		16'h16CA: out_word = 8'h5C;
		16'h16CB: out_word = 8'hE5;
		16'h16CC: out_word = 8'h21;
		16'h16CD: out_word = 8'h92;
		16'h16CE: out_word = 8'h5C;
		16'h16CF: out_word = 8'h22;
		16'h16D0: out_word = 8'h68;
		16'h16D1: out_word = 8'h5C;
		16'h16D2: out_word = 8'hE1;
		16'h16D3: out_word = 8'hC9;
		16'h16D4: out_word = 8'hED;
		16'h16D5: out_word = 8'h5B;
		16'h16D6: out_word = 8'h59;
		16'h16D7: out_word = 8'h5C;
		16'h16D8: out_word = 8'hC3;
		16'h16D9: out_word = 8'hE5;
		16'h16DA: out_word = 8'h19;
		16'h16DB: out_word = 8'h23;
		16'h16DC: out_word = 8'h7E;
		16'h16DD: out_word = 8'hA7;
		16'h16DE: out_word = 8'hC8;
		16'h16DF: out_word = 8'hB9;
		16'h16E0: out_word = 8'h23;
		16'h16E1: out_word = 8'h20;
		16'h16E2: out_word = 8'hF8;
		16'h16E3: out_word = 8'h37;
		16'h16E4: out_word = 8'hC9;
		16'h16E5: out_word = 8'hCD;
		16'h16E6: out_word = 8'h1E;
		16'h16E7: out_word = 8'h17;
		16'h16E8: out_word = 8'hCD;
		16'h16E9: out_word = 8'h01;
		16'h16EA: out_word = 8'h17;
		16'h16EB: out_word = 8'h01;
		16'h16EC: out_word = 8'h00;
		16'h16ED: out_word = 8'h00;
		16'h16EE: out_word = 8'h11;
		16'h16EF: out_word = 8'hE2;
		16'h16F0: out_word = 8'hA3;
		16'h16F1: out_word = 8'hEB;
		16'h16F2: out_word = 8'h19;
		16'h16F3: out_word = 8'h38;
		16'h16F4: out_word = 8'h07;
		16'h16F5: out_word = 8'h01;
		16'h16F6: out_word = 8'hD4;
		16'h16F7: out_word = 8'h15;
		16'h16F8: out_word = 8'h09;
		16'h16F9: out_word = 8'h4E;
		16'h16FA: out_word = 8'h23;
		16'h16FB: out_word = 8'h46;
		16'h16FC: out_word = 8'hEB;
		16'h16FD: out_word = 8'h71;
		16'h16FE: out_word = 8'h23;
		16'h16FF: out_word = 8'h70;
		16'h1700: out_word = 8'hC9;
		16'h1701: out_word = 8'hE5;
		16'h1702: out_word = 8'h2A;
		16'h1703: out_word = 8'h4F;
		16'h1704: out_word = 8'h5C;
		16'h1705: out_word = 8'h09;
		16'h1706: out_word = 8'h23;
		16'h1707: out_word = 8'h23;
		16'h1708: out_word = 8'h23;
		16'h1709: out_word = 8'h4E;
		16'h170A: out_word = 8'hEB;
		16'h170B: out_word = 8'h21;
		16'h170C: out_word = 8'h16;
		16'h170D: out_word = 8'h17;
		16'h170E: out_word = 8'hCD;
		16'h170F: out_word = 8'hDC;
		16'h1710: out_word = 8'h16;
		16'h1711: out_word = 8'h4E;
		16'h1712: out_word = 8'h06;
		16'h1713: out_word = 8'h00;
		16'h1714: out_word = 8'h09;
		16'h1715: out_word = 8'hE9;
		16'h1716: out_word = 8'h4B;
		16'h1717: out_word = 8'h05;
		16'h1718: out_word = 8'h53;
		16'h1719: out_word = 8'h03;
		16'h171A: out_word = 8'h50;
		16'h171B: out_word = 8'h01;
		16'h171C: out_word = 8'hE1;
		16'h171D: out_word = 8'hC9;
		16'h171E: out_word = 8'hCD;
		16'h171F: out_word = 8'h94;
		16'h1720: out_word = 8'h1E;
		16'h1721: out_word = 8'hFE;
		16'h1722: out_word = 8'h10;
		16'h1723: out_word = 8'h38;
		16'h1724: out_word = 8'h02;
		16'h1725: out_word = 8'hCF;
		16'h1726: out_word = 8'h17;
		16'h1727: out_word = 8'hC6;
		16'h1728: out_word = 8'h03;
		16'h1729: out_word = 8'h07;
		16'h172A: out_word = 8'h21;
		16'h172B: out_word = 8'h10;
		16'h172C: out_word = 8'h5C;
		16'h172D: out_word = 8'h4F;
		16'h172E: out_word = 8'h06;
		16'h172F: out_word = 8'h00;
		16'h1730: out_word = 8'h09;
		16'h1731: out_word = 8'h4E;
		16'h1732: out_word = 8'h23;
		16'h1733: out_word = 8'h46;
		16'h1734: out_word = 8'h2B;
		16'h1735: out_word = 8'hC9;
		16'h1736: out_word = 8'hEF;
		16'h1737: out_word = 8'h01;
		16'h1738: out_word = 8'h38;
		16'h1739: out_word = 8'hCD;
		16'h173A: out_word = 8'h1E;
		16'h173B: out_word = 8'h17;
		16'h173C: out_word = 8'h78;
		16'h173D: out_word = 8'hB1;
		16'h173E: out_word = 8'h28;
		16'h173F: out_word = 8'h16;
		16'h1740: out_word = 8'hEB;
		16'h1741: out_word = 8'h2A;
		16'h1742: out_word = 8'h4F;
		16'h1743: out_word = 8'h5C;
		16'h1744: out_word = 8'h09;
		16'h1745: out_word = 8'h23;
		16'h1746: out_word = 8'h23;
		16'h1747: out_word = 8'h23;
		16'h1748: out_word = 8'h7E;
		16'h1749: out_word = 8'hEB;
		16'h174A: out_word = 8'hFE;
		16'h174B: out_word = 8'h4B;
		16'h174C: out_word = 8'h28;
		16'h174D: out_word = 8'h08;
		16'h174E: out_word = 8'hFE;
		16'h174F: out_word = 8'h53;
		16'h1750: out_word = 8'h28;
		16'h1751: out_word = 8'h04;
		16'h1752: out_word = 8'hFE;
		16'h1753: out_word = 8'h50;
		16'h1754: out_word = 8'h20;
		16'h1755: out_word = 8'hCF;
		16'h1756: out_word = 8'hCD;
		16'h1757: out_word = 8'h5D;
		16'h1758: out_word = 8'h17;
		16'h1759: out_word = 8'h73;
		16'h175A: out_word = 8'h23;
		16'h175B: out_word = 8'h72;
		16'h175C: out_word = 8'hC9;
		16'h175D: out_word = 8'hE5;
		16'h175E: out_word = 8'hCD;
		16'h175F: out_word = 8'hF1;
		16'h1760: out_word = 8'h2B;
		16'h1761: out_word = 8'h78;
		16'h1762: out_word = 8'hB1;
		16'h1763: out_word = 8'h20;
		16'h1764: out_word = 8'h02;
		16'h1765: out_word = 8'hCF;
		16'h1766: out_word = 8'h0E;
		16'h1767: out_word = 8'hC5;
		16'h1768: out_word = 8'h1A;
		16'h1769: out_word = 8'hE6;
		16'h176A: out_word = 8'hDF;
		16'h176B: out_word = 8'h4F;
		16'h176C: out_word = 8'h21;
		16'h176D: out_word = 8'h7A;
		16'h176E: out_word = 8'h17;
		16'h176F: out_word = 8'hCD;
		16'h1770: out_word = 8'hDC;
		16'h1771: out_word = 8'h16;
		16'h1772: out_word = 8'h30;
		16'h1773: out_word = 8'hF1;
		16'h1774: out_word = 8'h4E;
		16'h1775: out_word = 8'h06;
		16'h1776: out_word = 8'h00;
		16'h1777: out_word = 8'h09;
		16'h1778: out_word = 8'hC1;
		16'h1779: out_word = 8'hE9;
		16'h177A: out_word = 8'h4B;
		16'h177B: out_word = 8'h06;
		16'h177C: out_word = 8'h53;
		16'h177D: out_word = 8'h08;
		16'h177E: out_word = 8'h50;
		16'h177F: out_word = 8'h0A;
		16'h1780: out_word = 8'h00;
		16'h1781: out_word = 8'h1E;
		16'h1782: out_word = 8'h01;
		16'h1783: out_word = 8'h18;
		16'h1784: out_word = 8'h06;
		16'h1785: out_word = 8'h1E;
		16'h1786: out_word = 8'h06;
		16'h1787: out_word = 8'h18;
		16'h1788: out_word = 8'h02;
		16'h1789: out_word = 8'h1E;
		16'h178A: out_word = 8'h10;
		16'h178B: out_word = 8'h0B;
		16'h178C: out_word = 8'h78;
		16'h178D: out_word = 8'hB1;
		16'h178E: out_word = 8'h20;
		16'h178F: out_word = 8'hD5;
		16'h1790: out_word = 8'h57;
		16'h1791: out_word = 8'hE1;
		16'h1792: out_word = 8'hC9;
		16'h1793: out_word = 8'h18;
		16'h1794: out_word = 8'h90;
		16'h1795: out_word = 8'hED;
		16'h1796: out_word = 8'h73;
		16'h1797: out_word = 8'h3F;
		16'h1798: out_word = 8'h5C;
		16'h1799: out_word = 8'hFD;
		16'h179A: out_word = 8'h36;
		16'h179B: out_word = 8'h02;
		16'h179C: out_word = 8'h10;
		16'h179D: out_word = 8'hCD;
		16'h179E: out_word = 8'hAF;
		16'h179F: out_word = 8'h0D;
		16'h17A0: out_word = 8'hFD;
		16'h17A1: out_word = 8'hCB;
		16'h17A2: out_word = 8'h02;
		16'h17A3: out_word = 8'hC6;
		16'h17A4: out_word = 8'hFD;
		16'h17A5: out_word = 8'h46;
		16'h17A6: out_word = 8'h31;
		16'h17A7: out_word = 8'hCD;
		16'h17A8: out_word = 8'h44;
		16'h17A9: out_word = 8'h0E;
		16'h17AA: out_word = 8'hFD;
		16'h17AB: out_word = 8'hCB;
		16'h17AC: out_word = 8'h02;
		16'h17AD: out_word = 8'h86;
		16'h17AE: out_word = 8'hFD;
		16'h17AF: out_word = 8'hCB;
		16'h17B0: out_word = 8'h30;
		16'h17B1: out_word = 8'hC6;
		16'h17B2: out_word = 8'h2A;
		16'h17B3: out_word = 8'h49;
		16'h17B4: out_word = 8'h5C;
		16'h17B5: out_word = 8'hED;
		16'h17B6: out_word = 8'h5B;
		16'h17B7: out_word = 8'h6C;
		16'h17B8: out_word = 8'h5C;
		16'h17B9: out_word = 8'hA7;
		16'h17BA: out_word = 8'hED;
		16'h17BB: out_word = 8'h52;
		16'h17BC: out_word = 8'h19;
		16'h17BD: out_word = 8'h38;
		16'h17BE: out_word = 8'h22;
		16'h17BF: out_word = 8'hD5;
		16'h17C0: out_word = 8'hCD;
		16'h17C1: out_word = 8'h6E;
		16'h17C2: out_word = 8'h19;
		16'h17C3: out_word = 8'h11;
		16'h17C4: out_word = 8'hC0;
		16'h17C5: out_word = 8'h02;
		16'h17C6: out_word = 8'hEB;
		16'h17C7: out_word = 8'hED;
		16'h17C8: out_word = 8'h52;
		16'h17C9: out_word = 8'hE3;
		16'h17CA: out_word = 8'hCD;
		16'h17CB: out_word = 8'h6E;
		16'h17CC: out_word = 8'h19;
		16'h17CD: out_word = 8'hC1;
		16'h17CE: out_word = 8'hC5;
		16'h17CF: out_word = 8'hCD;
		16'h17D0: out_word = 8'hB8;
		16'h17D1: out_word = 8'h19;
		16'h17D2: out_word = 8'hC1;
		16'h17D3: out_word = 8'h09;
		16'h17D4: out_word = 8'h38;
		16'h17D5: out_word = 8'h0E;
		16'h17D6: out_word = 8'hEB;
		16'h17D7: out_word = 8'h56;
		16'h17D8: out_word = 8'h23;
		16'h17D9: out_word = 8'h5E;
		16'h17DA: out_word = 8'h2B;
		16'h17DB: out_word = 8'hED;
		16'h17DC: out_word = 8'h53;
		16'h17DD: out_word = 8'h6C;
		16'h17DE: out_word = 8'h5C;
		16'h17DF: out_word = 8'h18;
		16'h17E0: out_word = 8'hED;
		16'h17E1: out_word = 8'h22;
		16'h17E2: out_word = 8'h6C;
		16'h17E3: out_word = 8'h5C;
		16'h17E4: out_word = 8'h2A;
		16'h17E5: out_word = 8'h6C;
		16'h17E6: out_word = 8'h5C;
		16'h17E7: out_word = 8'hCD;
		16'h17E8: out_word = 8'h6E;
		16'h17E9: out_word = 8'h19;
		16'h17EA: out_word = 8'h28;
		16'h17EB: out_word = 8'h01;
		16'h17EC: out_word = 8'hEB;
		16'h17ED: out_word = 8'hCD;
		16'h17EE: out_word = 8'h33;
		16'h17EF: out_word = 8'h18;
		16'h17F0: out_word = 8'hFD;
		16'h17F1: out_word = 8'hCB;
		16'h17F2: out_word = 8'h02;
		16'h17F3: out_word = 8'hA6;
		16'h17F4: out_word = 8'hC9;
		16'h17F5: out_word = 8'h3E;
		16'h17F6: out_word = 8'h03;
		16'h17F7: out_word = 8'h18;
		16'h17F8: out_word = 8'h02;
		16'h17F9: out_word = 8'h3E;
		16'h17FA: out_word = 8'h02;
		16'h17FB: out_word = 8'hFD;
		16'h17FC: out_word = 8'h36;
		16'h17FD: out_word = 8'h02;
		16'h17FE: out_word = 8'h00;
		16'h17FF: out_word = 8'hCD;
		16'h1800: out_word = 8'h30;
		16'h1801: out_word = 8'h25;
		16'h1802: out_word = 8'hC4;
		16'h1803: out_word = 8'h01;
		16'h1804: out_word = 8'h16;
		16'h1805: out_word = 8'hDF;
		16'h1806: out_word = 8'hCD;
		16'h1807: out_word = 8'h70;
		16'h1808: out_word = 8'h20;
		16'h1809: out_word = 8'h38;
		16'h180A: out_word = 8'h14;
		16'h180B: out_word = 8'hDF;
		16'h180C: out_word = 8'hFE;
		16'h180D: out_word = 8'h3B;
		16'h180E: out_word = 8'h28;
		16'h180F: out_word = 8'h04;
		16'h1810: out_word = 8'hFE;
		16'h1811: out_word = 8'h2C;
		16'h1812: out_word = 8'h20;
		16'h1813: out_word = 8'h06;
		16'h1814: out_word = 8'hE7;
		16'h1815: out_word = 8'hCD;
		16'h1816: out_word = 8'h82;
		16'h1817: out_word = 8'h1C;
		16'h1818: out_word = 8'h18;
		16'h1819: out_word = 8'h08;
		16'h181A: out_word = 8'hCD;
		16'h181B: out_word = 8'hE6;
		16'h181C: out_word = 8'h1C;
		16'h181D: out_word = 8'h18;
		16'h181E: out_word = 8'h03;
		16'h181F: out_word = 8'hCD;
		16'h1820: out_word = 8'hDE;
		16'h1821: out_word = 8'h1C;
		16'h1822: out_word = 8'hCD;
		16'h1823: out_word = 8'hEE;
		16'h1824: out_word = 8'h1B;
		16'h1825: out_word = 8'hCD;
		16'h1826: out_word = 8'h99;
		16'h1827: out_word = 8'h1E;
		16'h1828: out_word = 8'h78;
		16'h1829: out_word = 8'hE6;
		16'h182A: out_word = 8'h3F;
		16'h182B: out_word = 8'h67;
		16'h182C: out_word = 8'h69;
		16'h182D: out_word = 8'h22;
		16'h182E: out_word = 8'h49;
		16'h182F: out_word = 8'h5C;
		16'h1830: out_word = 8'hCD;
		16'h1831: out_word = 8'h6E;
		16'h1832: out_word = 8'h19;
		16'h1833: out_word = 8'h1E;
		16'h1834: out_word = 8'h01;
		16'h1835: out_word = 8'hCD;
		16'h1836: out_word = 8'h55;
		16'h1837: out_word = 8'h18;
		16'h1838: out_word = 8'hD7;
		16'h1839: out_word = 8'hFD;
		16'h183A: out_word = 8'hCB;
		16'h183B: out_word = 8'h02;
		16'h183C: out_word = 8'h66;
		16'h183D: out_word = 8'h28;
		16'h183E: out_word = 8'hF6;
		16'h183F: out_word = 8'h3A;
		16'h1840: out_word = 8'h6B;
		16'h1841: out_word = 8'h5C;
		16'h1842: out_word = 8'hFD;
		16'h1843: out_word = 8'h96;
		16'h1844: out_word = 8'h4F;
		16'h1845: out_word = 8'h20;
		16'h1846: out_word = 8'hEE;
		16'h1847: out_word = 8'hAB;
		16'h1848: out_word = 8'hC8;
		16'h1849: out_word = 8'hE5;
		16'h184A: out_word = 8'hD5;
		16'h184B: out_word = 8'h21;
		16'h184C: out_word = 8'h6C;
		16'h184D: out_word = 8'h5C;
		16'h184E: out_word = 8'hCD;
		16'h184F: out_word = 8'h0F;
		16'h1850: out_word = 8'h19;
		16'h1851: out_word = 8'hD1;
		16'h1852: out_word = 8'hE1;
		16'h1853: out_word = 8'h18;
		16'h1854: out_word = 8'hE0;
		16'h1855: out_word = 8'hED;
		16'h1856: out_word = 8'h4B;
		16'h1857: out_word = 8'h49;
		16'h1858: out_word = 8'h5C;
		16'h1859: out_word = 8'hCD;
		16'h185A: out_word = 8'h80;
		16'h185B: out_word = 8'h19;
		16'h185C: out_word = 8'h16;
		16'h185D: out_word = 8'h3E;
		16'h185E: out_word = 8'h28;
		16'h185F: out_word = 8'h05;
		16'h1860: out_word = 8'h11;
		16'h1861: out_word = 8'h00;
		16'h1862: out_word = 8'h00;
		16'h1863: out_word = 8'hCB;
		16'h1864: out_word = 8'h13;
		16'h1865: out_word = 8'hFD;
		16'h1866: out_word = 8'h73;
		16'h1867: out_word = 8'h2D;
		16'h1868: out_word = 8'h7E;
		16'h1869: out_word = 8'hFE;
		16'h186A: out_word = 8'h40;
		16'h186B: out_word = 8'hC1;
		16'h186C: out_word = 8'hD0;
		16'h186D: out_word = 8'hC5;
		16'h186E: out_word = 8'hCD;
		16'h186F: out_word = 8'h28;
		16'h1870: out_word = 8'h1A;
		16'h1871: out_word = 8'h23;
		16'h1872: out_word = 8'h23;
		16'h1873: out_word = 8'h23;
		16'h1874: out_word = 8'hFD;
		16'h1875: out_word = 8'hCB;
		16'h1876: out_word = 8'h01;
		16'h1877: out_word = 8'h86;
		16'h1878: out_word = 8'h7A;
		16'h1879: out_word = 8'hA7;
		16'h187A: out_word = 8'h28;
		16'h187B: out_word = 8'h05;
		16'h187C: out_word = 8'hD7;
		16'h187D: out_word = 8'hFD;
		16'h187E: out_word = 8'hCB;
		16'h187F: out_word = 8'h01;
		16'h1880: out_word = 8'hC6;
		16'h1881: out_word = 8'hD5;
		16'h1882: out_word = 8'hEB;
		16'h1883: out_word = 8'hFD;
		16'h1884: out_word = 8'hCB;
		16'h1885: out_word = 8'h30;
		16'h1886: out_word = 8'h96;
		16'h1887: out_word = 8'h21;
		16'h1888: out_word = 8'h3B;
		16'h1889: out_word = 8'h5C;
		16'h188A: out_word = 8'hCB;
		16'h188B: out_word = 8'h96;
		16'h188C: out_word = 8'hFD;
		16'h188D: out_word = 8'hCB;
		16'h188E: out_word = 8'h37;
		16'h188F: out_word = 8'h6E;
		16'h1890: out_word = 8'h28;
		16'h1891: out_word = 8'h02;
		16'h1892: out_word = 8'hCB;
		16'h1893: out_word = 8'hD6;
		16'h1894: out_word = 8'h2A;
		16'h1895: out_word = 8'h5F;
		16'h1896: out_word = 8'h5C;
		16'h1897: out_word = 8'hA7;
		16'h1898: out_word = 8'hED;
		16'h1899: out_word = 8'h52;
		16'h189A: out_word = 8'h20;
		16'h189B: out_word = 8'h05;
		16'h189C: out_word = 8'h3E;
		16'h189D: out_word = 8'h3F;
		16'h189E: out_word = 8'hCD;
		16'h189F: out_word = 8'hC1;
		16'h18A0: out_word = 8'h18;
		16'h18A1: out_word = 8'hCD;
		16'h18A2: out_word = 8'hE1;
		16'h18A3: out_word = 8'h18;
		16'h18A4: out_word = 8'hEB;
		16'h18A5: out_word = 8'h7E;
		16'h18A6: out_word = 8'hCD;
		16'h18A7: out_word = 8'hB6;
		16'h18A8: out_word = 8'h18;
		16'h18A9: out_word = 8'h23;
		16'h18AA: out_word = 8'hFE;
		16'h18AB: out_word = 8'h0D;
		16'h18AC: out_word = 8'h28;
		16'h18AD: out_word = 8'h06;
		16'h18AE: out_word = 8'hEB;
		16'h18AF: out_word = 8'hCD;
		16'h18B0: out_word = 8'h37;
		16'h18B1: out_word = 8'h19;
		16'h18B2: out_word = 8'h18;
		16'h18B3: out_word = 8'hE0;
		16'h18B4: out_word = 8'hD1;
		16'h18B5: out_word = 8'hC9;
		16'h18B6: out_word = 8'hFE;
		16'h18B7: out_word = 8'h0E;
		16'h18B8: out_word = 8'hC0;
		16'h18B9: out_word = 8'h23;
		16'h18BA: out_word = 8'h23;
		16'h18BB: out_word = 8'h23;
		16'h18BC: out_word = 8'h23;
		16'h18BD: out_word = 8'h23;
		16'h18BE: out_word = 8'h23;
		16'h18BF: out_word = 8'h7E;
		16'h18C0: out_word = 8'hC9;
		16'h18C1: out_word = 8'hD9;
		16'h18C2: out_word = 8'h2A;
		16'h18C3: out_word = 8'h8F;
		16'h18C4: out_word = 8'h5C;
		16'h18C5: out_word = 8'hE5;
		16'h18C6: out_word = 8'hCB;
		16'h18C7: out_word = 8'hBC;
		16'h18C8: out_word = 8'hCB;
		16'h18C9: out_word = 8'hFD;
		16'h18CA: out_word = 8'h22;
		16'h18CB: out_word = 8'h8F;
		16'h18CC: out_word = 8'h5C;
		16'h18CD: out_word = 8'h21;
		16'h18CE: out_word = 8'h91;
		16'h18CF: out_word = 8'h5C;
		16'h18D0: out_word = 8'h56;
		16'h18D1: out_word = 8'hD5;
		16'h18D2: out_word = 8'h36;
		16'h18D3: out_word = 8'h00;
		16'h18D4: out_word = 8'hCD;
		16'h18D5: out_word = 8'hF4;
		16'h18D6: out_word = 8'h09;
		16'h18D7: out_word = 8'hE1;
		16'h18D8: out_word = 8'hFD;
		16'h18D9: out_word = 8'h74;
		16'h18DA: out_word = 8'h57;
		16'h18DB: out_word = 8'hE1;
		16'h18DC: out_word = 8'h22;
		16'h18DD: out_word = 8'h8F;
		16'h18DE: out_word = 8'h5C;
		16'h18DF: out_word = 8'hD9;
		16'h18E0: out_word = 8'hC9;
		16'h18E1: out_word = 8'h2A;
		16'h18E2: out_word = 8'h5B;
		16'h18E3: out_word = 8'h5C;
		16'h18E4: out_word = 8'hA7;
		16'h18E5: out_word = 8'hED;
		16'h18E6: out_word = 8'h52;
		16'h18E7: out_word = 8'hC0;
		16'h18E8: out_word = 8'h3A;
		16'h18E9: out_word = 8'h41;
		16'h18EA: out_word = 8'h5C;
		16'h18EB: out_word = 8'hCB;
		16'h18EC: out_word = 8'h07;
		16'h18ED: out_word = 8'h28;
		16'h18EE: out_word = 8'h04;
		16'h18EF: out_word = 8'hC6;
		16'h18F0: out_word = 8'h43;
		16'h18F1: out_word = 8'h18;
		16'h18F2: out_word = 8'h16;
		16'h18F3: out_word = 8'h21;
		16'h18F4: out_word = 8'h3B;
		16'h18F5: out_word = 8'h5C;
		16'h18F6: out_word = 8'hCB;
		16'h18F7: out_word = 8'h9E;
		16'h18F8: out_word = 8'h3E;
		16'h18F9: out_word = 8'h4B;
		16'h18FA: out_word = 8'hCB;
		16'h18FB: out_word = 8'h56;
		16'h18FC: out_word = 8'h28;
		16'h18FD: out_word = 8'h0B;
		16'h18FE: out_word = 8'hCB;
		16'h18FF: out_word = 8'hDE;
		16'h1900: out_word = 8'h3C;
		16'h1901: out_word = 8'hFD;
		16'h1902: out_word = 8'hCB;
		16'h1903: out_word = 8'h30;
		16'h1904: out_word = 8'h5E;
		16'h1905: out_word = 8'h28;
		16'h1906: out_word = 8'h02;
		16'h1907: out_word = 8'h3E;
		16'h1908: out_word = 8'h43;
		16'h1909: out_word = 8'hD5;
		16'h190A: out_word = 8'hCD;
		16'h190B: out_word = 8'hC1;
		16'h190C: out_word = 8'h18;
		16'h190D: out_word = 8'hD1;
		16'h190E: out_word = 8'hC9;
		16'h190F: out_word = 8'h5E;
		16'h1910: out_word = 8'h23;
		16'h1911: out_word = 8'h56;
		16'h1912: out_word = 8'hE5;
		16'h1913: out_word = 8'hEB;
		16'h1914: out_word = 8'h23;
		16'h1915: out_word = 8'hCD;
		16'h1916: out_word = 8'h6E;
		16'h1917: out_word = 8'h19;
		16'h1918: out_word = 8'hCD;
		16'h1919: out_word = 8'h95;
		16'h191A: out_word = 8'h16;
		16'h191B: out_word = 8'hE1;
		16'h191C: out_word = 8'hFD;
		16'h191D: out_word = 8'hCB;
		16'h191E: out_word = 8'h37;
		16'h191F: out_word = 8'h6E;
		16'h1920: out_word = 8'hC0;
		16'h1921: out_word = 8'h72;
		16'h1922: out_word = 8'h2B;
		16'h1923: out_word = 8'h73;
		16'h1924: out_word = 8'hC9;
		16'h1925: out_word = 8'h7B;
		16'h1926: out_word = 8'hA7;
		16'h1927: out_word = 8'hF8;
		16'h1928: out_word = 8'h18;
		16'h1929: out_word = 8'h0D;
		16'h192A: out_word = 8'hAF;
		16'h192B: out_word = 8'h09;
		16'h192C: out_word = 8'h3C;
		16'h192D: out_word = 8'h38;
		16'h192E: out_word = 8'hFC;
		16'h192F: out_word = 8'hED;
		16'h1930: out_word = 8'h42;
		16'h1931: out_word = 8'h3D;
		16'h1932: out_word = 8'h28;
		16'h1933: out_word = 8'hF1;
		16'h1934: out_word = 8'hC3;
		16'h1935: out_word = 8'hEF;
		16'h1936: out_word = 8'h15;
		16'h1937: out_word = 8'hCD;
		16'h1938: out_word = 8'h1B;
		16'h1939: out_word = 8'h2D;
		16'h193A: out_word = 8'h30;
		16'h193B: out_word = 8'h30;
		16'h193C: out_word = 8'hFE;
		16'h193D: out_word = 8'h21;
		16'h193E: out_word = 8'h38;
		16'h193F: out_word = 8'h2C;
		16'h1940: out_word = 8'hFD;
		16'h1941: out_word = 8'hCB;
		16'h1942: out_word = 8'h01;
		16'h1943: out_word = 8'h96;
		16'h1944: out_word = 8'hFE;
		16'h1945: out_word = 8'hCB;
		16'h1946: out_word = 8'h28;
		16'h1947: out_word = 8'h24;
		16'h1948: out_word = 8'hFE;
		16'h1949: out_word = 8'h3A;
		16'h194A: out_word = 8'h20;
		16'h194B: out_word = 8'h0E;
		16'h194C: out_word = 8'hFD;
		16'h194D: out_word = 8'hCB;
		16'h194E: out_word = 8'h37;
		16'h194F: out_word = 8'h6E;
		16'h1950: out_word = 8'h20;
		16'h1951: out_word = 8'h16;
		16'h1952: out_word = 8'hFD;
		16'h1953: out_word = 8'hCB;
		16'h1954: out_word = 8'h30;
		16'h1955: out_word = 8'h56;
		16'h1956: out_word = 8'h28;
		16'h1957: out_word = 8'h14;
		16'h1958: out_word = 8'h18;
		16'h1959: out_word = 8'h0E;
		16'h195A: out_word = 8'hFE;
		16'h195B: out_word = 8'h22;
		16'h195C: out_word = 8'h20;
		16'h195D: out_word = 8'h0A;
		16'h195E: out_word = 8'hF5;
		16'h195F: out_word = 8'h3A;
		16'h1960: out_word = 8'h6A;
		16'h1961: out_word = 8'h5C;
		16'h1962: out_word = 8'hEE;
		16'h1963: out_word = 8'h04;
		16'h1964: out_word = 8'h32;
		16'h1965: out_word = 8'h6A;
		16'h1966: out_word = 8'h5C;
		16'h1967: out_word = 8'hF1;
		16'h1968: out_word = 8'hFD;
		16'h1969: out_word = 8'hCB;
		16'h196A: out_word = 8'h01;
		16'h196B: out_word = 8'hD6;
		16'h196C: out_word = 8'hD7;
		16'h196D: out_word = 8'hC9;
		16'h196E: out_word = 8'hE5;
		16'h196F: out_word = 8'h2A;
		16'h1970: out_word = 8'h53;
		16'h1971: out_word = 8'h5C;
		16'h1972: out_word = 8'h54;
		16'h1973: out_word = 8'h5D;
		16'h1974: out_word = 8'hC1;
		16'h1975: out_word = 8'hCD;
		16'h1976: out_word = 8'h80;
		16'h1977: out_word = 8'h19;
		16'h1978: out_word = 8'hD0;
		16'h1979: out_word = 8'hC5;
		16'h197A: out_word = 8'hCD;
		16'h197B: out_word = 8'hB8;
		16'h197C: out_word = 8'h19;
		16'h197D: out_word = 8'hEB;
		16'h197E: out_word = 8'h18;
		16'h197F: out_word = 8'hF4;
		16'h1980: out_word = 8'h7E;
		16'h1981: out_word = 8'hB8;
		16'h1982: out_word = 8'hC0;
		16'h1983: out_word = 8'h23;
		16'h1984: out_word = 8'h7E;
		16'h1985: out_word = 8'h2B;
		16'h1986: out_word = 8'hB9;
		16'h1987: out_word = 8'hC9;
		16'h1988: out_word = 8'h23;
		16'h1989: out_word = 8'h23;
		16'h198A: out_word = 8'h23;
		16'h198B: out_word = 8'h22;
		16'h198C: out_word = 8'h5D;
		16'h198D: out_word = 8'h5C;
		16'h198E: out_word = 8'h0E;
		16'h198F: out_word = 8'h00;
		16'h1990: out_word = 8'h15;
		16'h1991: out_word = 8'hC8;
		16'h1992: out_word = 8'hE7;
		16'h1993: out_word = 8'hBB;
		16'h1994: out_word = 8'h20;
		16'h1995: out_word = 8'h04;
		16'h1996: out_word = 8'hA7;
		16'h1997: out_word = 8'hC9;
		16'h1998: out_word = 8'h23;
		16'h1999: out_word = 8'h7E;
		16'h199A: out_word = 8'hCD;
		16'h199B: out_word = 8'hB6;
		16'h199C: out_word = 8'h18;
		16'h199D: out_word = 8'h22;
		16'h199E: out_word = 8'h5D;
		16'h199F: out_word = 8'h5C;
		16'h19A0: out_word = 8'hFE;
		16'h19A1: out_word = 8'h22;
		16'h19A2: out_word = 8'h20;
		16'h19A3: out_word = 8'h01;
		16'h19A4: out_word = 8'h0D;
		16'h19A5: out_word = 8'hFE;
		16'h19A6: out_word = 8'h3A;
		16'h19A7: out_word = 8'h28;
		16'h19A8: out_word = 8'h04;
		16'h19A9: out_word = 8'hFE;
		16'h19AA: out_word = 8'hCB;
		16'h19AB: out_word = 8'h20;
		16'h19AC: out_word = 8'h04;
		16'h19AD: out_word = 8'hCB;
		16'h19AE: out_word = 8'h41;
		16'h19AF: out_word = 8'h28;
		16'h19B0: out_word = 8'hDF;
		16'h19B1: out_word = 8'hFE;
		16'h19B2: out_word = 8'h0D;
		16'h19B3: out_word = 8'h20;
		16'h19B4: out_word = 8'hE3;
		16'h19B5: out_word = 8'h15;
		16'h19B6: out_word = 8'h37;
		16'h19B7: out_word = 8'hC9;
		16'h19B8: out_word = 8'hE5;
		16'h19B9: out_word = 8'h7E;
		16'h19BA: out_word = 8'hFE;
		16'h19BB: out_word = 8'h40;
		16'h19BC: out_word = 8'h38;
		16'h19BD: out_word = 8'h17;
		16'h19BE: out_word = 8'hCB;
		16'h19BF: out_word = 8'h6F;
		16'h19C0: out_word = 8'h28;
		16'h19C1: out_word = 8'h14;
		16'h19C2: out_word = 8'h87;
		16'h19C3: out_word = 8'hFA;
		16'h19C4: out_word = 8'hC7;
		16'h19C5: out_word = 8'h19;
		16'h19C6: out_word = 8'h3F;
		16'h19C7: out_word = 8'h01;
		16'h19C8: out_word = 8'h05;
		16'h19C9: out_word = 8'h00;
		16'h19CA: out_word = 8'h30;
		16'h19CB: out_word = 8'h02;
		16'h19CC: out_word = 8'h0E;
		16'h19CD: out_word = 8'h12;
		16'h19CE: out_word = 8'h17;
		16'h19CF: out_word = 8'h23;
		16'h19D0: out_word = 8'h7E;
		16'h19D1: out_word = 8'h30;
		16'h19D2: out_word = 8'hFB;
		16'h19D3: out_word = 8'h18;
		16'h19D4: out_word = 8'h06;
		16'h19D5: out_word = 8'h23;
		16'h19D6: out_word = 8'h23;
		16'h19D7: out_word = 8'h4E;
		16'h19D8: out_word = 8'h23;
		16'h19D9: out_word = 8'h46;
		16'h19DA: out_word = 8'h23;
		16'h19DB: out_word = 8'h09;
		16'h19DC: out_word = 8'hD1;
		16'h19DD: out_word = 8'hA7;
		16'h19DE: out_word = 8'hED;
		16'h19DF: out_word = 8'h52;
		16'h19E0: out_word = 8'h44;
		16'h19E1: out_word = 8'h4D;
		16'h19E2: out_word = 8'h19;
		16'h19E3: out_word = 8'hEB;
		16'h19E4: out_word = 8'hC9;
		16'h19E5: out_word = 8'hCD;
		16'h19E6: out_word = 8'hDD;
		16'h19E7: out_word = 8'h19;
		16'h19E8: out_word = 8'hC5;
		16'h19E9: out_word = 8'h78;
		16'h19EA: out_word = 8'h2F;
		16'h19EB: out_word = 8'h47;
		16'h19EC: out_word = 8'h79;
		16'h19ED: out_word = 8'h2F;
		16'h19EE: out_word = 8'h4F;
		16'h19EF: out_word = 8'h03;
		16'h19F0: out_word = 8'hCD;
		16'h19F1: out_word = 8'h64;
		16'h19F2: out_word = 8'h16;
		16'h19F3: out_word = 8'hEB;
		16'h19F4: out_word = 8'hE1;
		16'h19F5: out_word = 8'h19;
		16'h19F6: out_word = 8'hD5;
		16'h19F7: out_word = 8'hED;
		16'h19F8: out_word = 8'hB0;
		16'h19F9: out_word = 8'hE1;
		16'h19FA: out_word = 8'hC9;
		16'h19FB: out_word = 8'h2A;
		16'h19FC: out_word = 8'h59;
		16'h19FD: out_word = 8'h5C;
		16'h19FE: out_word = 8'h2B;
		16'h19FF: out_word = 8'h22;
		16'h1A00: out_word = 8'h5D;
		16'h1A01: out_word = 8'h5C;
		16'h1A02: out_word = 8'hE7;
		16'h1A03: out_word = 8'h21;
		16'h1A04: out_word = 8'h92;
		16'h1A05: out_word = 8'h5C;
		16'h1A06: out_word = 8'h22;
		16'h1A07: out_word = 8'h65;
		16'h1A08: out_word = 8'h5C;
		16'h1A09: out_word = 8'hCD;
		16'h1A0A: out_word = 8'h3B;
		16'h1A0B: out_word = 8'h2D;
		16'h1A0C: out_word = 8'hCD;
		16'h1A0D: out_word = 8'hA2;
		16'h1A0E: out_word = 8'h2D;
		16'h1A0F: out_word = 8'h38;
		16'h1A10: out_word = 8'h04;
		16'h1A11: out_word = 8'h21;
		16'h1A12: out_word = 8'hF0;
		16'h1A13: out_word = 8'hD8;
		16'h1A14: out_word = 8'h09;
		16'h1A15: out_word = 8'hDA;
		16'h1A16: out_word = 8'h8A;
		16'h1A17: out_word = 8'h1C;
		16'h1A18: out_word = 8'hC3;
		16'h1A19: out_word = 8'hC5;
		16'h1A1A: out_word = 8'h16;
		16'h1A1B: out_word = 8'hD5;
		16'h1A1C: out_word = 8'hE5;
		16'h1A1D: out_word = 8'hAF;
		16'h1A1E: out_word = 8'hCB;
		16'h1A1F: out_word = 8'h78;
		16'h1A20: out_word = 8'h20;
		16'h1A21: out_word = 8'h20;
		16'h1A22: out_word = 8'h60;
		16'h1A23: out_word = 8'h69;
		16'h1A24: out_word = 8'h1E;
		16'h1A25: out_word = 8'hFF;
		16'h1A26: out_word = 8'h18;
		16'h1A27: out_word = 8'h08;
		16'h1A28: out_word = 8'hD5;
		16'h1A29: out_word = 8'h56;
		16'h1A2A: out_word = 8'h23;
		16'h1A2B: out_word = 8'h5E;
		16'h1A2C: out_word = 8'hE5;
		16'h1A2D: out_word = 8'hEB;
		16'h1A2E: out_word = 8'h1E;
		16'h1A2F: out_word = 8'h20;
		16'h1A30: out_word = 8'h01;
		16'h1A31: out_word = 8'h18;
		16'h1A32: out_word = 8'hFC;
		16'h1A33: out_word = 8'hCD;
		16'h1A34: out_word = 8'h2A;
		16'h1A35: out_word = 8'h19;
		16'h1A36: out_word = 8'h01;
		16'h1A37: out_word = 8'h9C;
		16'h1A38: out_word = 8'hFF;
		16'h1A39: out_word = 8'hCD;
		16'h1A3A: out_word = 8'h2A;
		16'h1A3B: out_word = 8'h19;
		16'h1A3C: out_word = 8'h0E;
		16'h1A3D: out_word = 8'hF6;
		16'h1A3E: out_word = 8'hCD;
		16'h1A3F: out_word = 8'h2A;
		16'h1A40: out_word = 8'h19;
		16'h1A41: out_word = 8'h7D;
		16'h1A42: out_word = 8'hCD;
		16'h1A43: out_word = 8'hEF;
		16'h1A44: out_word = 8'h15;
		16'h1A45: out_word = 8'hE1;
		16'h1A46: out_word = 8'hD1;
		16'h1A47: out_word = 8'hC9;
		16'h1A48: out_word = 8'hB1;
		16'h1A49: out_word = 8'hCB;
		16'h1A4A: out_word = 8'hBC;
		16'h1A4B: out_word = 8'hBF;
		16'h1A4C: out_word = 8'hC4;
		16'h1A4D: out_word = 8'hAF;
		16'h1A4E: out_word = 8'hB4;
		16'h1A4F: out_word = 8'h93;
		16'h1A50: out_word = 8'h91;
		16'h1A51: out_word = 8'h92;
		16'h1A52: out_word = 8'h95;
		16'h1A53: out_word = 8'h98;
		16'h1A54: out_word = 8'h98;
		16'h1A55: out_word = 8'h98;
		16'h1A56: out_word = 8'h98;
		16'h1A57: out_word = 8'h98;
		16'h1A58: out_word = 8'h98;
		16'h1A59: out_word = 8'h98;
		16'h1A5A: out_word = 8'h7F;
		16'h1A5B: out_word = 8'h81;
		16'h1A5C: out_word = 8'h2E;
		16'h1A5D: out_word = 8'h6C;
		16'h1A5E: out_word = 8'h6E;
		16'h1A5F: out_word = 8'h70;
		16'h1A60: out_word = 8'h48;
		16'h1A61: out_word = 8'h94;
		16'h1A62: out_word = 8'h56;
		16'h1A63: out_word = 8'h3F;
		16'h1A64: out_word = 8'h41;
		16'h1A65: out_word = 8'h2B;
		16'h1A66: out_word = 8'h17;
		16'h1A67: out_word = 8'h1F;
		16'h1A68: out_word = 8'h37;
		16'h1A69: out_word = 8'h77;
		16'h1A6A: out_word = 8'h44;
		16'h1A6B: out_word = 8'h0F;
		16'h1A6C: out_word = 8'h59;
		16'h1A6D: out_word = 8'h2B;
		16'h1A6E: out_word = 8'h43;
		16'h1A6F: out_word = 8'h2D;
		16'h1A70: out_word = 8'h51;
		16'h1A71: out_word = 8'h3A;
		16'h1A72: out_word = 8'h6D;
		16'h1A73: out_word = 8'h42;
		16'h1A74: out_word = 8'h0D;
		16'h1A75: out_word = 8'h49;
		16'h1A76: out_word = 8'h5C;
		16'h1A77: out_word = 8'h44;
		16'h1A78: out_word = 8'h15;
		16'h1A79: out_word = 8'h5D;
		16'h1A7A: out_word = 8'h01;
		16'h1A7B: out_word = 8'h3D;
		16'h1A7C: out_word = 8'h02;
		16'h1A7D: out_word = 8'h06;
		16'h1A7E: out_word = 8'h00;
		16'h1A7F: out_word = 8'h67;
		16'h1A80: out_word = 8'h1E;
		16'h1A81: out_word = 8'h06;
		16'h1A82: out_word = 8'hCB;
		16'h1A83: out_word = 8'h05;
		16'h1A84: out_word = 8'hF0;
		16'h1A85: out_word = 8'h1C;
		16'h1A86: out_word = 8'h06;
		16'h1A87: out_word = 8'h00;
		16'h1A88: out_word = 8'hED;
		16'h1A89: out_word = 8'h1E;
		16'h1A8A: out_word = 8'h00;
		16'h1A8B: out_word = 8'hEE;
		16'h1A8C: out_word = 8'h1C;
		16'h1A8D: out_word = 8'h00;
		16'h1A8E: out_word = 8'h23;
		16'h1A8F: out_word = 8'h1F;
		16'h1A90: out_word = 8'h04;
		16'h1A91: out_word = 8'h3D;
		16'h1A92: out_word = 8'h06;
		16'h1A93: out_word = 8'hCC;
		16'h1A94: out_word = 8'h06;
		16'h1A95: out_word = 8'h05;
		16'h1A96: out_word = 8'h03;
		16'h1A97: out_word = 8'h1D;
		16'h1A98: out_word = 8'h04;
		16'h1A99: out_word = 8'h00;
		16'h1A9A: out_word = 8'hAB;
		16'h1A9B: out_word = 8'h1D;
		16'h1A9C: out_word = 8'h05;
		16'h1A9D: out_word = 8'hCD;
		16'h1A9E: out_word = 8'h1F;
		16'h1A9F: out_word = 8'h05;
		16'h1AA0: out_word = 8'h89;
		16'h1AA1: out_word = 8'h20;
		16'h1AA2: out_word = 8'h05;
		16'h1AA3: out_word = 8'h02;
		16'h1AA4: out_word = 8'h2C;
		16'h1AA5: out_word = 8'h05;
		16'h1AA6: out_word = 8'hB2;
		16'h1AA7: out_word = 8'h1B;
		16'h1AA8: out_word = 8'h00;
		16'h1AA9: out_word = 8'hB7;
		16'h1AAA: out_word = 8'h11;
		16'h1AAB: out_word = 8'h03;
		16'h1AAC: out_word = 8'hA1;
		16'h1AAD: out_word = 8'h1E;
		16'h1AAE: out_word = 8'h05;
		16'h1AAF: out_word = 8'hF9;
		16'h1AB0: out_word = 8'h17;
		16'h1AB1: out_word = 8'h08;
		16'h1AB2: out_word = 8'h00;
		16'h1AB3: out_word = 8'h80;
		16'h1AB4: out_word = 8'h1E;
		16'h1AB5: out_word = 8'h03;
		16'h1AB6: out_word = 8'h4F;
		16'h1AB7: out_word = 8'h1E;
		16'h1AB8: out_word = 8'h00;
		16'h1AB9: out_word = 8'h5F;
		16'h1ABA: out_word = 8'h1E;
		16'h1ABB: out_word = 8'h03;
		16'h1ABC: out_word = 8'hAC;
		16'h1ABD: out_word = 8'h1E;
		16'h1ABE: out_word = 8'h00;
		16'h1ABF: out_word = 8'h6B;
		16'h1AC0: out_word = 8'h0D;
		16'h1AC1: out_word = 8'h09;
		16'h1AC2: out_word = 8'h00;
		16'h1AC3: out_word = 8'hDC;
		16'h1AC4: out_word = 8'h22;
		16'h1AC5: out_word = 8'h06;
		16'h1AC6: out_word = 8'h00;
		16'h1AC7: out_word = 8'h3A;
		16'h1AC8: out_word = 8'h1F;
		16'h1AC9: out_word = 8'h05;
		16'h1ACA: out_word = 8'hED;
		16'h1ACB: out_word = 8'h1D;
		16'h1ACC: out_word = 8'h05;
		16'h1ACD: out_word = 8'h27;
		16'h1ACE: out_word = 8'h1E;
		16'h1ACF: out_word = 8'h03;
		16'h1AD0: out_word = 8'h42;
		16'h1AD1: out_word = 8'h1E;
		16'h1AD2: out_word = 8'h09;
		16'h1AD3: out_word = 8'h05;
		16'h1AD4: out_word = 8'h82;
		16'h1AD5: out_word = 8'h23;
		16'h1AD6: out_word = 8'h00;
		16'h1AD7: out_word = 8'hAC;
		16'h1AD8: out_word = 8'h0E;
		16'h1AD9: out_word = 8'h05;
		16'h1ADA: out_word = 8'hC9;
		16'h1ADB: out_word = 8'h1F;
		16'h1ADC: out_word = 8'h05;
		16'h1ADD: out_word = 8'hF5;
		16'h1ADE: out_word = 8'h17;
		16'h1ADF: out_word = 8'h0B;
		16'h1AE0: out_word = 8'h0B;
		16'h1AE1: out_word = 8'h0B;
		16'h1AE2: out_word = 8'h0B;
		16'h1AE3: out_word = 8'h08;
		16'h1AE4: out_word = 8'h00;
		16'h1AE5: out_word = 8'hF8;
		16'h1AE6: out_word = 8'h03;
		16'h1AE7: out_word = 8'h09;
		16'h1AE8: out_word = 8'h05;
		16'h1AE9: out_word = 8'h20;
		16'h1AEA: out_word = 8'h23;
		16'h1AEB: out_word = 8'h07;
		16'h1AEC: out_word = 8'h07;
		16'h1AED: out_word = 8'h07;
		16'h1AEE: out_word = 8'h07;
		16'h1AEF: out_word = 8'h07;
		16'h1AF0: out_word = 8'h07;
		16'h1AF1: out_word = 8'h08;
		16'h1AF2: out_word = 8'h00;
		16'h1AF3: out_word = 8'h7A;
		16'h1AF4: out_word = 8'h1E;
		16'h1AF5: out_word = 8'h06;
		16'h1AF6: out_word = 8'h00;
		16'h1AF7: out_word = 8'h94;
		16'h1AF8: out_word = 8'h22;
		16'h1AF9: out_word = 8'h05;
		16'h1AFA: out_word = 8'h60;
		16'h1AFB: out_word = 8'h1F;
		16'h1AFC: out_word = 8'h06;
		16'h1AFD: out_word = 8'h2C;
		16'h1AFE: out_word = 8'h0A;
		16'h1AFF: out_word = 8'h00;
		16'h1B00: out_word = 8'h36;
		16'h1B01: out_word = 8'h17;
		16'h1B02: out_word = 8'h06;
		16'h1B03: out_word = 8'h00;
		16'h1B04: out_word = 8'hE5;
		16'h1B05: out_word = 8'h16;
		16'h1B06: out_word = 8'h0A;
		16'h1B07: out_word = 8'h00;
		16'h1B08: out_word = 8'h93;
		16'h1B09: out_word = 8'h17;
		16'h1B0A: out_word = 8'h0A;
		16'h1B0B: out_word = 8'h2C;
		16'h1B0C: out_word = 8'h0A;
		16'h1B0D: out_word = 8'h00;
		16'h1B0E: out_word = 8'h93;
		16'h1B0F: out_word = 8'h17;
		16'h1B10: out_word = 8'h0A;
		16'h1B11: out_word = 8'h00;
		16'h1B12: out_word = 8'h93;
		16'h1B13: out_word = 8'h17;
		16'h1B14: out_word = 8'h00;
		16'h1B15: out_word = 8'h93;
		16'h1B16: out_word = 8'h17;
		16'h1B17: out_word = 8'hFD;
		16'h1B18: out_word = 8'hCB;
		16'h1B19: out_word = 8'h01;
		16'h1B1A: out_word = 8'hBE;
		16'h1B1B: out_word = 8'hCD;
		16'h1B1C: out_word = 8'hFB;
		16'h1B1D: out_word = 8'h19;
		16'h1B1E: out_word = 8'hAF;
		16'h1B1F: out_word = 8'h32;
		16'h1B20: out_word = 8'h47;
		16'h1B21: out_word = 8'h5C;
		16'h1B22: out_word = 8'h3D;
		16'h1B23: out_word = 8'h32;
		16'h1B24: out_word = 8'h3A;
		16'h1B25: out_word = 8'h5C;
		16'h1B26: out_word = 8'h18;
		16'h1B27: out_word = 8'h01;
		16'h1B28: out_word = 8'hE7;
		16'h1B29: out_word = 8'hCD;
		16'h1B2A: out_word = 8'hBF;
		16'h1B2B: out_word = 8'h16;
		16'h1B2C: out_word = 8'hFD;
		16'h1B2D: out_word = 8'h34;
		16'h1B2E: out_word = 8'h0D;
		16'h1B2F: out_word = 8'hFA;
		16'h1B30: out_word = 8'h8A;
		16'h1B31: out_word = 8'h1C;
		16'h1B32: out_word = 8'hDF;
		16'h1B33: out_word = 8'h06;
		16'h1B34: out_word = 8'h00;
		16'h1B35: out_word = 8'hFE;
		16'h1B36: out_word = 8'h0D;
		16'h1B37: out_word = 8'h28;
		16'h1B38: out_word = 8'h7A;
		16'h1B39: out_word = 8'hFE;
		16'h1B3A: out_word = 8'h3A;
		16'h1B3B: out_word = 8'h28;
		16'h1B3C: out_word = 8'hEB;
		16'h1B3D: out_word = 8'h21;
		16'h1B3E: out_word = 8'h76;
		16'h1B3F: out_word = 8'h1B;
		16'h1B40: out_word = 8'hE5;
		16'h1B41: out_word = 8'h4F;
		16'h1B42: out_word = 8'hE7;
		16'h1B43: out_word = 8'h79;
		16'h1B44: out_word = 8'hD6;
		16'h1B45: out_word = 8'hCE;
		16'h1B46: out_word = 8'hDA;
		16'h1B47: out_word = 8'h8A;
		16'h1B48: out_word = 8'h1C;
		16'h1B49: out_word = 8'h4F;
		16'h1B4A: out_word = 8'h21;
		16'h1B4B: out_word = 8'h48;
		16'h1B4C: out_word = 8'h1A;
		16'h1B4D: out_word = 8'h09;
		16'h1B4E: out_word = 8'h4E;
		16'h1B4F: out_word = 8'h09;
		16'h1B50: out_word = 8'h18;
		16'h1B51: out_word = 8'h03;
		16'h1B52: out_word = 8'h2A;
		16'h1B53: out_word = 8'h74;
		16'h1B54: out_word = 8'h5C;
		16'h1B55: out_word = 8'h7E;
		16'h1B56: out_word = 8'h23;
		16'h1B57: out_word = 8'h22;
		16'h1B58: out_word = 8'h74;
		16'h1B59: out_word = 8'h5C;
		16'h1B5A: out_word = 8'h01;
		16'h1B5B: out_word = 8'h52;
		16'h1B5C: out_word = 8'h1B;
		16'h1B5D: out_word = 8'hC5;
		16'h1B5E: out_word = 8'h4F;
		16'h1B5F: out_word = 8'hFE;
		16'h1B60: out_word = 8'h20;
		16'h1B61: out_word = 8'h30;
		16'h1B62: out_word = 8'h0C;
		16'h1B63: out_word = 8'h21;
		16'h1B64: out_word = 8'h01;
		16'h1B65: out_word = 8'h1C;
		16'h1B66: out_word = 8'h06;
		16'h1B67: out_word = 8'h00;
		16'h1B68: out_word = 8'h09;
		16'h1B69: out_word = 8'h4E;
		16'h1B6A: out_word = 8'h09;
		16'h1B6B: out_word = 8'hE5;
		16'h1B6C: out_word = 8'hDF;
		16'h1B6D: out_word = 8'h05;
		16'h1B6E: out_word = 8'hC9;
		16'h1B6F: out_word = 8'hDF;
		16'h1B70: out_word = 8'hB9;
		16'h1B71: out_word = 8'hC2;
		16'h1B72: out_word = 8'h8A;
		16'h1B73: out_word = 8'h1C;
		16'h1B74: out_word = 8'hE7;
		16'h1B75: out_word = 8'hC9;
		16'h1B76: out_word = 8'hCD;
		16'h1B77: out_word = 8'h54;
		16'h1B78: out_word = 8'h1F;
		16'h1B79: out_word = 8'h38;
		16'h1B7A: out_word = 8'h02;
		16'h1B7B: out_word = 8'hCF;
		16'h1B7C: out_word = 8'h14;
		16'h1B7D: out_word = 8'hCD;
		16'h1B7E: out_word = 8'h4D;
		16'h1B7F: out_word = 8'h3B;
		16'h1B80: out_word = 8'h00;
		16'h1B81: out_word = 8'h20;
		16'h1B82: out_word = 8'h71;
		16'h1B83: out_word = 8'h2A;
		16'h1B84: out_word = 8'h42;
		16'h1B85: out_word = 8'h5C;
		16'h1B86: out_word = 8'hCB;
		16'h1B87: out_word = 8'h7C;
		16'h1B88: out_word = 8'h28;
		16'h1B89: out_word = 8'h14;
		16'h1B8A: out_word = 8'h21;
		16'h1B8B: out_word = 8'hFE;
		16'h1B8C: out_word = 8'hFF;
		16'h1B8D: out_word = 8'h22;
		16'h1B8E: out_word = 8'h45;
		16'h1B8F: out_word = 8'h5C;
		16'h1B90: out_word = 8'h2A;
		16'h1B91: out_word = 8'h61;
		16'h1B92: out_word = 8'h5C;
		16'h1B93: out_word = 8'h2B;
		16'h1B94: out_word = 8'hED;
		16'h1B95: out_word = 8'h5B;
		16'h1B96: out_word = 8'h59;
		16'h1B97: out_word = 8'h5C;
		16'h1B98: out_word = 8'h1B;
		16'h1B99: out_word = 8'h3A;
		16'h1B9A: out_word = 8'h44;
		16'h1B9B: out_word = 8'h5C;
		16'h1B9C: out_word = 8'h18;
		16'h1B9D: out_word = 8'h33;
		16'h1B9E: out_word = 8'hCD;
		16'h1B9F: out_word = 8'h6E;
		16'h1BA0: out_word = 8'h19;
		16'h1BA1: out_word = 8'h3A;
		16'h1BA2: out_word = 8'h44;
		16'h1BA3: out_word = 8'h5C;
		16'h1BA4: out_word = 8'h28;
		16'h1BA5: out_word = 8'h19;
		16'h1BA6: out_word = 8'hA7;
		16'h1BA7: out_word = 8'h20;
		16'h1BA8: out_word = 8'h43;
		16'h1BA9: out_word = 8'h47;
		16'h1BAA: out_word = 8'h7E;
		16'h1BAB: out_word = 8'hE6;
		16'h1BAC: out_word = 8'hC0;
		16'h1BAD: out_word = 8'h78;
		16'h1BAE: out_word = 8'h28;
		16'h1BAF: out_word = 8'h0F;
		16'h1BB0: out_word = 8'hCF;
		16'h1BB1: out_word = 8'hFF;
		16'h1BB2: out_word = 8'hC1;
		16'h1BB3: out_word = 8'hCD;
		16'h1BB4: out_word = 8'h30;
		16'h1BB5: out_word = 8'h25;
		16'h1BB6: out_word = 8'hC8;
		16'h1BB7: out_word = 8'h2A;
		16'h1BB8: out_word = 8'h55;
		16'h1BB9: out_word = 8'h5C;
		16'h1BBA: out_word = 8'h3E;
		16'h1BBB: out_word = 8'hC0;
		16'h1BBC: out_word = 8'hA6;
		16'h1BBD: out_word = 8'hC0;
		16'h1BBE: out_word = 8'hAF;
		16'h1BBF: out_word = 8'hFE;
		16'h1BC0: out_word = 8'h01;
		16'h1BC1: out_word = 8'hCE;
		16'h1BC2: out_word = 8'h00;
		16'h1BC3: out_word = 8'h56;
		16'h1BC4: out_word = 8'h23;
		16'h1BC5: out_word = 8'h5E;
		16'h1BC6: out_word = 8'hED;
		16'h1BC7: out_word = 8'h53;
		16'h1BC8: out_word = 8'h45;
		16'h1BC9: out_word = 8'h5C;
		16'h1BCA: out_word = 8'h23;
		16'h1BCB: out_word = 8'h5E;
		16'h1BCC: out_word = 8'h23;
		16'h1BCD: out_word = 8'h56;
		16'h1BCE: out_word = 8'hEB;
		16'h1BCF: out_word = 8'h19;
		16'h1BD0: out_word = 8'h23;
		16'h1BD1: out_word = 8'h22;
		16'h1BD2: out_word = 8'h55;
		16'h1BD3: out_word = 8'h5C;
		16'h1BD4: out_word = 8'hEB;
		16'h1BD5: out_word = 8'h22;
		16'h1BD6: out_word = 8'h5D;
		16'h1BD7: out_word = 8'h5C;
		16'h1BD8: out_word = 8'h57;
		16'h1BD9: out_word = 8'h1E;
		16'h1BDA: out_word = 8'h00;
		16'h1BDB: out_word = 8'hFD;
		16'h1BDC: out_word = 8'h36;
		16'h1BDD: out_word = 8'h0A;
		16'h1BDE: out_word = 8'hFF;
		16'h1BDF: out_word = 8'h15;
		16'h1BE0: out_word = 8'hFD;
		16'h1BE1: out_word = 8'h72;
		16'h1BE2: out_word = 8'h0D;
		16'h1BE3: out_word = 8'hCA;
		16'h1BE4: out_word = 8'h28;
		16'h1BE5: out_word = 8'h1B;
		16'h1BE6: out_word = 8'h14;
		16'h1BE7: out_word = 8'hCD;
		16'h1BE8: out_word = 8'h8B;
		16'h1BE9: out_word = 8'h19;
		16'h1BEA: out_word = 8'h28;
		16'h1BEB: out_word = 8'h08;
		16'h1BEC: out_word = 8'hCF;
		16'h1BED: out_word = 8'h16;
		16'h1BEE: out_word = 8'hCD;
		16'h1BEF: out_word = 8'h30;
		16'h1BF0: out_word = 8'h25;
		16'h1BF1: out_word = 8'hC0;
		16'h1BF2: out_word = 8'hC1;
		16'h1BF3: out_word = 8'hC1;
		16'h1BF4: out_word = 8'hCD;
		16'h1BF5: out_word = 8'h5D;
		16'h1BF6: out_word = 8'h3B;
		16'h1BF7: out_word = 8'h28;
		16'h1BF8: out_word = 8'hBA;
		16'h1BF9: out_word = 8'hFE;
		16'h1BFA: out_word = 8'h3A;
		16'h1BFB: out_word = 8'hCA;
		16'h1BFC: out_word = 8'h28;
		16'h1BFD: out_word = 8'h1B;
		16'h1BFE: out_word = 8'hC3;
		16'h1BFF: out_word = 8'h8A;
		16'h1C00: out_word = 8'h1C;
		16'h1C01: out_word = 8'h0F;
		16'h1C02: out_word = 8'h1D;
		16'h1C03: out_word = 8'h4B;
		16'h1C04: out_word = 8'h09;
		16'h1C05: out_word = 8'h67;
		16'h1C06: out_word = 8'h0B;
		16'h1C07: out_word = 8'h7B;
		16'h1C08: out_word = 8'h8E;
		16'h1C09: out_word = 8'h71;
		16'h1C0A: out_word = 8'hB4;
		16'h1C0B: out_word = 8'h81;
		16'h1C0C: out_word = 8'hCF;
		16'h1C0D: out_word = 8'hCD;
		16'h1C0E: out_word = 8'hDE;
		16'h1C0F: out_word = 8'h1C;
		16'h1C10: out_word = 8'hBF;
		16'h1C11: out_word = 8'hC1;
		16'h1C12: out_word = 8'hCC;
		16'h1C13: out_word = 8'hEE;
		16'h1C14: out_word = 8'h1B;
		16'h1C15: out_word = 8'hEB;
		16'h1C16: out_word = 8'h2A;
		16'h1C17: out_word = 8'h74;
		16'h1C18: out_word = 8'h5C;
		16'h1C19: out_word = 8'h4E;
		16'h1C1A: out_word = 8'h23;
		16'h1C1B: out_word = 8'h46;
		16'h1C1C: out_word = 8'hEB;
		16'h1C1D: out_word = 8'hC5;
		16'h1C1E: out_word = 8'hC9;
		16'h1C1F: out_word = 8'hCD;
		16'h1C20: out_word = 8'hB2;
		16'h1C21: out_word = 8'h28;
		16'h1C22: out_word = 8'hFD;
		16'h1C23: out_word = 8'h36;
		16'h1C24: out_word = 8'h37;
		16'h1C25: out_word = 8'h00;
		16'h1C26: out_word = 8'h30;
		16'h1C27: out_word = 8'h08;
		16'h1C28: out_word = 8'hFD;
		16'h1C29: out_word = 8'hCB;
		16'h1C2A: out_word = 8'h37;
		16'h1C2B: out_word = 8'hCE;
		16'h1C2C: out_word = 8'h20;
		16'h1C2D: out_word = 8'h18;
		16'h1C2E: out_word = 8'hCF;
		16'h1C2F: out_word = 8'h01;
		16'h1C30: out_word = 8'hCC;
		16'h1C31: out_word = 8'h96;
		16'h1C32: out_word = 8'h29;
		16'h1C33: out_word = 8'hFD;
		16'h1C34: out_word = 8'hCB;
		16'h1C35: out_word = 8'h01;
		16'h1C36: out_word = 8'h76;
		16'h1C37: out_word = 8'h20;
		16'h1C38: out_word = 8'h0D;
		16'h1C39: out_word = 8'hAF;
		16'h1C3A: out_word = 8'hCD;
		16'h1C3B: out_word = 8'h30;
		16'h1C3C: out_word = 8'h25;
		16'h1C3D: out_word = 8'hC4;
		16'h1C3E: out_word = 8'hF1;
		16'h1C3F: out_word = 8'h2B;
		16'h1C40: out_word = 8'h21;
		16'h1C41: out_word = 8'h71;
		16'h1C42: out_word = 8'h5C;
		16'h1C43: out_word = 8'hB6;
		16'h1C44: out_word = 8'h77;
		16'h1C45: out_word = 8'hEB;
		16'h1C46: out_word = 8'hED;
		16'h1C47: out_word = 8'h43;
		16'h1C48: out_word = 8'h72;
		16'h1C49: out_word = 8'h5C;
		16'h1C4A: out_word = 8'h22;
		16'h1C4B: out_word = 8'h4D;
		16'h1C4C: out_word = 8'h5C;
		16'h1C4D: out_word = 8'hC9;
		16'h1C4E: out_word = 8'hC1;
		16'h1C4F: out_word = 8'hCD;
		16'h1C50: out_word = 8'h56;
		16'h1C51: out_word = 8'h1C;
		16'h1C52: out_word = 8'hCD;
		16'h1C53: out_word = 8'hEE;
		16'h1C54: out_word = 8'h1B;
		16'h1C55: out_word = 8'hC9;
		16'h1C56: out_word = 8'h3A;
		16'h1C57: out_word = 8'h3B;
		16'h1C58: out_word = 8'h5C;
		16'h1C59: out_word = 8'hF5;
		16'h1C5A: out_word = 8'hCD;
		16'h1C5B: out_word = 8'hFB;
		16'h1C5C: out_word = 8'h24;
		16'h1C5D: out_word = 8'hF1;
		16'h1C5E: out_word = 8'hFD;
		16'h1C5F: out_word = 8'h56;
		16'h1C60: out_word = 8'h01;
		16'h1C61: out_word = 8'hAA;
		16'h1C62: out_word = 8'hE6;
		16'h1C63: out_word = 8'h40;
		16'h1C64: out_word = 8'h20;
		16'h1C65: out_word = 8'h24;
		16'h1C66: out_word = 8'hCB;
		16'h1C67: out_word = 8'h7A;
		16'h1C68: out_word = 8'hC2;
		16'h1C69: out_word = 8'hFF;
		16'h1C6A: out_word = 8'h2A;
		16'h1C6B: out_word = 8'hC9;
		16'h1C6C: out_word = 8'hCD;
		16'h1C6D: out_word = 8'hB2;
		16'h1C6E: out_word = 8'h28;
		16'h1C6F: out_word = 8'hF5;
		16'h1C70: out_word = 8'h79;
		16'h1C71: out_word = 8'hF6;
		16'h1C72: out_word = 8'h9F;
		16'h1C73: out_word = 8'h3C;
		16'h1C74: out_word = 8'h20;
		16'h1C75: out_word = 8'h14;
		16'h1C76: out_word = 8'hF1;
		16'h1C77: out_word = 8'h18;
		16'h1C78: out_word = 8'hA9;
		16'h1C79: out_word = 8'hE7;
		16'h1C7A: out_word = 8'hCD;
		16'h1C7B: out_word = 8'h82;
		16'h1C7C: out_word = 8'h1C;
		16'h1C7D: out_word = 8'hFE;
		16'h1C7E: out_word = 8'h2C;
		16'h1C7F: out_word = 8'h20;
		16'h1C80: out_word = 8'h09;
		16'h1C81: out_word = 8'hE7;
		16'h1C82: out_word = 8'hCD;
		16'h1C83: out_word = 8'hFB;
		16'h1C84: out_word = 8'h24;
		16'h1C85: out_word = 8'hFD;
		16'h1C86: out_word = 8'hCB;
		16'h1C87: out_word = 8'h01;
		16'h1C88: out_word = 8'h76;
		16'h1C89: out_word = 8'hC0;
		16'h1C8A: out_word = 8'hCF;
		16'h1C8B: out_word = 8'h0B;
		16'h1C8C: out_word = 8'hCD;
		16'h1C8D: out_word = 8'hFB;
		16'h1C8E: out_word = 8'h24;
		16'h1C8F: out_word = 8'hFD;
		16'h1C90: out_word = 8'hCB;
		16'h1C91: out_word = 8'h01;
		16'h1C92: out_word = 8'h76;
		16'h1C93: out_word = 8'hC8;
		16'h1C94: out_word = 8'h18;
		16'h1C95: out_word = 8'hF4;
		16'h1C96: out_word = 8'hFD;
		16'h1C97: out_word = 8'hCB;
		16'h1C98: out_word = 8'h01;
		16'h1C99: out_word = 8'h7E;
		16'h1C9A: out_word = 8'hFD;
		16'h1C9B: out_word = 8'hCB;
		16'h1C9C: out_word = 8'h02;
		16'h1C9D: out_word = 8'h86;
		16'h1C9E: out_word = 8'hC4;
		16'h1C9F: out_word = 8'h4D;
		16'h1CA0: out_word = 8'h0D;
		16'h1CA1: out_word = 8'hF1;
		16'h1CA2: out_word = 8'h3A;
		16'h1CA3: out_word = 8'h74;
		16'h1CA4: out_word = 8'h5C;
		16'h1CA5: out_word = 8'hD6;
		16'h1CA6: out_word = 8'h13;
		16'h1CA7: out_word = 8'hCD;
		16'h1CA8: out_word = 8'hFC;
		16'h1CA9: out_word = 8'h21;
		16'h1CAA: out_word = 8'hCD;
		16'h1CAB: out_word = 8'hEE;
		16'h1CAC: out_word = 8'h1B;
		16'h1CAD: out_word = 8'h2A;
		16'h1CAE: out_word = 8'h8F;
		16'h1CAF: out_word = 8'h5C;
		16'h1CB0: out_word = 8'h22;
		16'h1CB1: out_word = 8'h8D;
		16'h1CB2: out_word = 8'h5C;
		16'h1CB3: out_word = 8'h21;
		16'h1CB4: out_word = 8'h91;
		16'h1CB5: out_word = 8'h5C;
		16'h1CB6: out_word = 8'h7E;
		16'h1CB7: out_word = 8'h07;
		16'h1CB8: out_word = 8'hAE;
		16'h1CB9: out_word = 8'hE6;
		16'h1CBA: out_word = 8'hAA;
		16'h1CBB: out_word = 8'hAE;
		16'h1CBC: out_word = 8'h77;
		16'h1CBD: out_word = 8'hC9;
		16'h1CBE: out_word = 8'hCD;
		16'h1CBF: out_word = 8'h30;
		16'h1CC0: out_word = 8'h25;
		16'h1CC1: out_word = 8'h28;
		16'h1CC2: out_word = 8'h13;
		16'h1CC3: out_word = 8'hFD;
		16'h1CC4: out_word = 8'hCB;
		16'h1CC5: out_word = 8'h02;
		16'h1CC6: out_word = 8'h86;
		16'h1CC7: out_word = 8'hCD;
		16'h1CC8: out_word = 8'h4D;
		16'h1CC9: out_word = 8'h0D;
		16'h1CCA: out_word = 8'h21;
		16'h1CCB: out_word = 8'h90;
		16'h1CCC: out_word = 8'h5C;
		16'h1CCD: out_word = 8'h7E;
		16'h1CCE: out_word = 8'hF6;
		16'h1CCF: out_word = 8'hF8;
		16'h1CD0: out_word = 8'h77;
		16'h1CD1: out_word = 8'hFD;
		16'h1CD2: out_word = 8'hCB;
		16'h1CD3: out_word = 8'h57;
		16'h1CD4: out_word = 8'hB6;
		16'h1CD5: out_word = 8'hDF;
		16'h1CD6: out_word = 8'hCD;
		16'h1CD7: out_word = 8'hE2;
		16'h1CD8: out_word = 8'h21;
		16'h1CD9: out_word = 8'h18;
		16'h1CDA: out_word = 8'h9F;
		16'h1CDB: out_word = 8'hC3;
		16'h1CDC: out_word = 8'h05;
		16'h1CDD: out_word = 8'h06;
		16'h1CDE: out_word = 8'hFE;
		16'h1CDF: out_word = 8'h0D;
		16'h1CE0: out_word = 8'h28;
		16'h1CE1: out_word = 8'h04;
		16'h1CE2: out_word = 8'hFE;
		16'h1CE3: out_word = 8'h3A;
		16'h1CE4: out_word = 8'h20;
		16'h1CE5: out_word = 8'h9C;
		16'h1CE6: out_word = 8'hCD;
		16'h1CE7: out_word = 8'h30;
		16'h1CE8: out_word = 8'h25;
		16'h1CE9: out_word = 8'hC8;
		16'h1CEA: out_word = 8'hEF;
		16'h1CEB: out_word = 8'hA0;
		16'h1CEC: out_word = 8'h38;
		16'h1CED: out_word = 8'hC9;
		16'h1CEE: out_word = 8'hCF;
		16'h1CEF: out_word = 8'h08;
		16'h1CF0: out_word = 8'hC1;
		16'h1CF1: out_word = 8'hCD;
		16'h1CF2: out_word = 8'h30;
		16'h1CF3: out_word = 8'h25;
		16'h1CF4: out_word = 8'h28;
		16'h1CF5: out_word = 8'h0A;
		16'h1CF6: out_word = 8'hEF;
		16'h1CF7: out_word = 8'h02;
		16'h1CF8: out_word = 8'h38;
		16'h1CF9: out_word = 8'hEB;
		16'h1CFA: out_word = 8'hCD;
		16'h1CFB: out_word = 8'hE9;
		16'h1CFC: out_word = 8'h34;
		16'h1CFD: out_word = 8'hDA;
		16'h1CFE: out_word = 8'hB3;
		16'h1CFF: out_word = 8'h1B;
		16'h1D00: out_word = 8'hC3;
		16'h1D01: out_word = 8'h29;
		16'h1D02: out_word = 8'h1B;
		16'h1D03: out_word = 8'hFE;
		16'h1D04: out_word = 8'hCD;
		16'h1D05: out_word = 8'h20;
		16'h1D06: out_word = 8'h09;
		16'h1D07: out_word = 8'hE7;
		16'h1D08: out_word = 8'hCD;
		16'h1D09: out_word = 8'h82;
		16'h1D0A: out_word = 8'h1C;
		16'h1D0B: out_word = 8'hCD;
		16'h1D0C: out_word = 8'hEE;
		16'h1D0D: out_word = 8'h1B;
		16'h1D0E: out_word = 8'h18;
		16'h1D0F: out_word = 8'h06;
		16'h1D10: out_word = 8'hCD;
		16'h1D11: out_word = 8'hEE;
		16'h1D12: out_word = 8'h1B;
		16'h1D13: out_word = 8'hEF;
		16'h1D14: out_word = 8'hA1;
		16'h1D15: out_word = 8'h38;
		16'h1D16: out_word = 8'hEF;
		16'h1D17: out_word = 8'hC0;
		16'h1D18: out_word = 8'h02;
		16'h1D19: out_word = 8'h01;
		16'h1D1A: out_word = 8'hE0;
		16'h1D1B: out_word = 8'h01;
		16'h1D1C: out_word = 8'h38;
		16'h1D1D: out_word = 8'hCD;
		16'h1D1E: out_word = 8'hFF;
		16'h1D1F: out_word = 8'h2A;
		16'h1D20: out_word = 8'h22;
		16'h1D21: out_word = 8'h68;
		16'h1D22: out_word = 8'h5C;
		16'h1D23: out_word = 8'h2B;
		16'h1D24: out_word = 8'h7E;
		16'h1D25: out_word = 8'hCB;
		16'h1D26: out_word = 8'hFE;
		16'h1D27: out_word = 8'h01;
		16'h1D28: out_word = 8'h06;
		16'h1D29: out_word = 8'h00;
		16'h1D2A: out_word = 8'h09;
		16'h1D2B: out_word = 8'h07;
		16'h1D2C: out_word = 8'h38;
		16'h1D2D: out_word = 8'h06;
		16'h1D2E: out_word = 8'h0E;
		16'h1D2F: out_word = 8'h0D;
		16'h1D30: out_word = 8'hCD;
		16'h1D31: out_word = 8'h55;
		16'h1D32: out_word = 8'h16;
		16'h1D33: out_word = 8'h23;
		16'h1D34: out_word = 8'hE5;
		16'h1D35: out_word = 8'hEF;
		16'h1D36: out_word = 8'h02;
		16'h1D37: out_word = 8'h02;
		16'h1D38: out_word = 8'h38;
		16'h1D39: out_word = 8'hE1;
		16'h1D3A: out_word = 8'hEB;
		16'h1D3B: out_word = 8'h0E;
		16'h1D3C: out_word = 8'h0A;
		16'h1D3D: out_word = 8'hED;
		16'h1D3E: out_word = 8'hB0;
		16'h1D3F: out_word = 8'h2A;
		16'h1D40: out_word = 8'h45;
		16'h1D41: out_word = 8'h5C;
		16'h1D42: out_word = 8'hEB;
		16'h1D43: out_word = 8'h73;
		16'h1D44: out_word = 8'h23;
		16'h1D45: out_word = 8'h72;
		16'h1D46: out_word = 8'hFD;
		16'h1D47: out_word = 8'h56;
		16'h1D48: out_word = 8'h0D;
		16'h1D49: out_word = 8'h14;
		16'h1D4A: out_word = 8'h23;
		16'h1D4B: out_word = 8'h72;
		16'h1D4C: out_word = 8'hCD;
		16'h1D4D: out_word = 8'hDA;
		16'h1D4E: out_word = 8'h1D;
		16'h1D4F: out_word = 8'hD0;
		16'h1D50: out_word = 8'hFD;
		16'h1D51: out_word = 8'h46;
		16'h1D52: out_word = 8'h38;
		16'h1D53: out_word = 8'h2A;
		16'h1D54: out_word = 8'h45;
		16'h1D55: out_word = 8'h5C;
		16'h1D56: out_word = 8'h22;
		16'h1D57: out_word = 8'h42;
		16'h1D58: out_word = 8'h5C;
		16'h1D59: out_word = 8'h3A;
		16'h1D5A: out_word = 8'h47;
		16'h1D5B: out_word = 8'h5C;
		16'h1D5C: out_word = 8'hED;
		16'h1D5D: out_word = 8'h44;
		16'h1D5E: out_word = 8'h57;
		16'h1D5F: out_word = 8'h2A;
		16'h1D60: out_word = 8'h5D;
		16'h1D61: out_word = 8'h5C;
		16'h1D62: out_word = 8'h1E;
		16'h1D63: out_word = 8'hF3;
		16'h1D64: out_word = 8'hC5;
		16'h1D65: out_word = 8'hED;
		16'h1D66: out_word = 8'h4B;
		16'h1D67: out_word = 8'h55;
		16'h1D68: out_word = 8'h5C;
		16'h1D69: out_word = 8'hCD;
		16'h1D6A: out_word = 8'h86;
		16'h1D6B: out_word = 8'h1D;
		16'h1D6C: out_word = 8'hED;
		16'h1D6D: out_word = 8'h43;
		16'h1D6E: out_word = 8'h55;
		16'h1D6F: out_word = 8'h5C;
		16'h1D70: out_word = 8'hC1;
		16'h1D71: out_word = 8'h38;
		16'h1D72: out_word = 8'h11;
		16'h1D73: out_word = 8'hE7;
		16'h1D74: out_word = 8'hF6;
		16'h1D75: out_word = 8'h20;
		16'h1D76: out_word = 8'hB8;
		16'h1D77: out_word = 8'h28;
		16'h1D78: out_word = 8'h03;
		16'h1D79: out_word = 8'hE7;
		16'h1D7A: out_word = 8'h18;
		16'h1D7B: out_word = 8'hE8;
		16'h1D7C: out_word = 8'hE7;
		16'h1D7D: out_word = 8'h3E;
		16'h1D7E: out_word = 8'h01;
		16'h1D7F: out_word = 8'h92;
		16'h1D80: out_word = 8'h32;
		16'h1D81: out_word = 8'h44;
		16'h1D82: out_word = 8'h5C;
		16'h1D83: out_word = 8'hC9;
		16'h1D84: out_word = 8'hCF;
		16'h1D85: out_word = 8'h11;
		16'h1D86: out_word = 8'h7E;
		16'h1D87: out_word = 8'hFE;
		16'h1D88: out_word = 8'h3A;
		16'h1D89: out_word = 8'h28;
		16'h1D8A: out_word = 8'h18;
		16'h1D8B: out_word = 8'h23;
		16'h1D8C: out_word = 8'h7E;
		16'h1D8D: out_word = 8'hE6;
		16'h1D8E: out_word = 8'hC0;
		16'h1D8F: out_word = 8'h37;
		16'h1D90: out_word = 8'hC0;
		16'h1D91: out_word = 8'h46;
		16'h1D92: out_word = 8'h23;
		16'h1D93: out_word = 8'h4E;
		16'h1D94: out_word = 8'hED;
		16'h1D95: out_word = 8'h43;
		16'h1D96: out_word = 8'h42;
		16'h1D97: out_word = 8'h5C;
		16'h1D98: out_word = 8'h23;
		16'h1D99: out_word = 8'h4E;
		16'h1D9A: out_word = 8'h23;
		16'h1D9B: out_word = 8'h46;
		16'h1D9C: out_word = 8'hE5;
		16'h1D9D: out_word = 8'h09;
		16'h1D9E: out_word = 8'h44;
		16'h1D9F: out_word = 8'h4D;
		16'h1DA0: out_word = 8'hE1;
		16'h1DA1: out_word = 8'h16;
		16'h1DA2: out_word = 8'h00;
		16'h1DA3: out_word = 8'hC5;
		16'h1DA4: out_word = 8'hCD;
		16'h1DA5: out_word = 8'h8B;
		16'h1DA6: out_word = 8'h19;
		16'h1DA7: out_word = 8'hC1;
		16'h1DA8: out_word = 8'hD0;
		16'h1DA9: out_word = 8'h18;
		16'h1DAA: out_word = 8'hE0;
		16'h1DAB: out_word = 8'hFD;
		16'h1DAC: out_word = 8'hCB;
		16'h1DAD: out_word = 8'h37;
		16'h1DAE: out_word = 8'h4E;
		16'h1DAF: out_word = 8'hC2;
		16'h1DB0: out_word = 8'h2E;
		16'h1DB1: out_word = 8'h1C;
		16'h1DB2: out_word = 8'h2A;
		16'h1DB3: out_word = 8'h4D;
		16'h1DB4: out_word = 8'h5C;
		16'h1DB5: out_word = 8'hCB;
		16'h1DB6: out_word = 8'h7E;
		16'h1DB7: out_word = 8'h28;
		16'h1DB8: out_word = 8'h1F;
		16'h1DB9: out_word = 8'h23;
		16'h1DBA: out_word = 8'h22;
		16'h1DBB: out_word = 8'h68;
		16'h1DBC: out_word = 8'h5C;
		16'h1DBD: out_word = 8'hEF;
		16'h1DBE: out_word = 8'hE0;
		16'h1DBF: out_word = 8'hE2;
		16'h1DC0: out_word = 8'h0F;
		16'h1DC1: out_word = 8'hC0;
		16'h1DC2: out_word = 8'h02;
		16'h1DC3: out_word = 8'h38;
		16'h1DC4: out_word = 8'hCD;
		16'h1DC5: out_word = 8'hDA;
		16'h1DC6: out_word = 8'h1D;
		16'h1DC7: out_word = 8'hD8;
		16'h1DC8: out_word = 8'h2A;
		16'h1DC9: out_word = 8'h68;
		16'h1DCA: out_word = 8'h5C;
		16'h1DCB: out_word = 8'h11;
		16'h1DCC: out_word = 8'h0F;
		16'h1DCD: out_word = 8'h00;
		16'h1DCE: out_word = 8'h19;
		16'h1DCF: out_word = 8'h5E;
		16'h1DD0: out_word = 8'h23;
		16'h1DD1: out_word = 8'h56;
		16'h1DD2: out_word = 8'h23;
		16'h1DD3: out_word = 8'h66;
		16'h1DD4: out_word = 8'hEB;
		16'h1DD5: out_word = 8'hC3;
		16'h1DD6: out_word = 8'h73;
		16'h1DD7: out_word = 8'h1E;
		16'h1DD8: out_word = 8'hCF;
		16'h1DD9: out_word = 8'h00;
		16'h1DDA: out_word = 8'hEF;
		16'h1DDB: out_word = 8'hE1;
		16'h1DDC: out_word = 8'hE0;
		16'h1DDD: out_word = 8'hE2;
		16'h1DDE: out_word = 8'h36;
		16'h1DDF: out_word = 8'h00;
		16'h1DE0: out_word = 8'h02;
		16'h1DE1: out_word = 8'h01;
		16'h1DE2: out_word = 8'h03;
		16'h1DE3: out_word = 8'h37;
		16'h1DE4: out_word = 8'h00;
		16'h1DE5: out_word = 8'h04;
		16'h1DE6: out_word = 8'h38;
		16'h1DE7: out_word = 8'hA7;
		16'h1DE8: out_word = 8'hC9;
		16'h1DE9: out_word = 8'h38;
		16'h1DEA: out_word = 8'h37;
		16'h1DEB: out_word = 8'hC9;
		16'h1DEC: out_word = 8'hE7;
		16'h1DED: out_word = 8'hCD;
		16'h1DEE: out_word = 8'h1F;
		16'h1DEF: out_word = 8'h1C;
		16'h1DF0: out_word = 8'hCD;
		16'h1DF1: out_word = 8'h30;
		16'h1DF2: out_word = 8'h25;
		16'h1DF3: out_word = 8'h28;
		16'h1DF4: out_word = 8'h29;
		16'h1DF5: out_word = 8'hDF;
		16'h1DF6: out_word = 8'h22;
		16'h1DF7: out_word = 8'h5F;
		16'h1DF8: out_word = 8'h5C;
		16'h1DF9: out_word = 8'h2A;
		16'h1DFA: out_word = 8'h57;
		16'h1DFB: out_word = 8'h5C;
		16'h1DFC: out_word = 8'h7E;
		16'h1DFD: out_word = 8'hFE;
		16'h1DFE: out_word = 8'h2C;
		16'h1DFF: out_word = 8'h28;
		16'h1E00: out_word = 8'h09;
		16'h1E01: out_word = 8'h1E;
		16'h1E02: out_word = 8'hE4;
		16'h1E03: out_word = 8'hCD;
		16'h1E04: out_word = 8'h86;
		16'h1E05: out_word = 8'h1D;
		16'h1E06: out_word = 8'h30;
		16'h1E07: out_word = 8'h02;
		16'h1E08: out_word = 8'hCF;
		16'h1E09: out_word = 8'h0D;
		16'h1E0A: out_word = 8'hCD;
		16'h1E0B: out_word = 8'h77;
		16'h1E0C: out_word = 8'h00;
		16'h1E0D: out_word = 8'hCD;
		16'h1E0E: out_word = 8'h56;
		16'h1E0F: out_word = 8'h1C;
		16'h1E10: out_word = 8'hDF;
		16'h1E11: out_word = 8'h22;
		16'h1E12: out_word = 8'h57;
		16'h1E13: out_word = 8'h5C;
		16'h1E14: out_word = 8'h2A;
		16'h1E15: out_word = 8'h5F;
		16'h1E16: out_word = 8'h5C;
		16'h1E17: out_word = 8'hFD;
		16'h1E18: out_word = 8'h36;
		16'h1E19: out_word = 8'h26;
		16'h1E1A: out_word = 8'h00;
		16'h1E1B: out_word = 8'hCD;
		16'h1E1C: out_word = 8'h78;
		16'h1E1D: out_word = 8'h00;
		16'h1E1E: out_word = 8'hDF;
		16'h1E1F: out_word = 8'hFE;
		16'h1E20: out_word = 8'h2C;
		16'h1E21: out_word = 8'h28;
		16'h1E22: out_word = 8'hC9;
		16'h1E23: out_word = 8'hCD;
		16'h1E24: out_word = 8'hEE;
		16'h1E25: out_word = 8'h1B;
		16'h1E26: out_word = 8'hC9;
		16'h1E27: out_word = 8'hCD;
		16'h1E28: out_word = 8'h30;
		16'h1E29: out_word = 8'h25;
		16'h1E2A: out_word = 8'h20;
		16'h1E2B: out_word = 8'h0B;
		16'h1E2C: out_word = 8'hCD;
		16'h1E2D: out_word = 8'hFB;
		16'h1E2E: out_word = 8'h24;
		16'h1E2F: out_word = 8'hFE;
		16'h1E30: out_word = 8'h2C;
		16'h1E31: out_word = 8'hC4;
		16'h1E32: out_word = 8'hEE;
		16'h1E33: out_word = 8'h1B;
		16'h1E34: out_word = 8'hE7;
		16'h1E35: out_word = 8'h18;
		16'h1E36: out_word = 8'hF5;
		16'h1E37: out_word = 8'h3E;
		16'h1E38: out_word = 8'hE4;
		16'h1E39: out_word = 8'h47;
		16'h1E3A: out_word = 8'hED;
		16'h1E3B: out_word = 8'hB9;
		16'h1E3C: out_word = 8'h11;
		16'h1E3D: out_word = 8'h00;
		16'h1E3E: out_word = 8'h02;
		16'h1E3F: out_word = 8'hC3;
		16'h1E40: out_word = 8'h8B;
		16'h1E41: out_word = 8'h19;
		16'h1E42: out_word = 8'hCD;
		16'h1E43: out_word = 8'h99;
		16'h1E44: out_word = 8'h1E;
		16'h1E45: out_word = 8'h60;
		16'h1E46: out_word = 8'h69;
		16'h1E47: out_word = 8'hCD;
		16'h1E48: out_word = 8'h6E;
		16'h1E49: out_word = 8'h19;
		16'h1E4A: out_word = 8'h2B;
		16'h1E4B: out_word = 8'h22;
		16'h1E4C: out_word = 8'h57;
		16'h1E4D: out_word = 8'h5C;
		16'h1E4E: out_word = 8'hC9;
		16'h1E4F: out_word = 8'hCD;
		16'h1E50: out_word = 8'h99;
		16'h1E51: out_word = 8'h1E;
		16'h1E52: out_word = 8'h78;
		16'h1E53: out_word = 8'hB1;
		16'h1E54: out_word = 8'h20;
		16'h1E55: out_word = 8'h04;
		16'h1E56: out_word = 8'hED;
		16'h1E57: out_word = 8'h4B;
		16'h1E58: out_word = 8'h78;
		16'h1E59: out_word = 8'h5C;
		16'h1E5A: out_word = 8'hED;
		16'h1E5B: out_word = 8'h43;
		16'h1E5C: out_word = 8'h76;
		16'h1E5D: out_word = 8'h5C;
		16'h1E5E: out_word = 8'hC9;
		16'h1E5F: out_word = 8'h2A;
		16'h1E60: out_word = 8'h6E;
		16'h1E61: out_word = 8'h5C;
		16'h1E62: out_word = 8'hFD;
		16'h1E63: out_word = 8'h56;
		16'h1E64: out_word = 8'h36;
		16'h1E65: out_word = 8'h18;
		16'h1E66: out_word = 8'h0C;
		16'h1E67: out_word = 8'hCD;
		16'h1E68: out_word = 8'h99;
		16'h1E69: out_word = 8'h1E;
		16'h1E6A: out_word = 8'h60;
		16'h1E6B: out_word = 8'h69;
		16'h1E6C: out_word = 8'h16;
		16'h1E6D: out_word = 8'h00;
		16'h1E6E: out_word = 8'h7C;
		16'h1E6F: out_word = 8'hFE;
		16'h1E70: out_word = 8'hF0;
		16'h1E71: out_word = 8'h30;
		16'h1E72: out_word = 8'h2C;
		16'h1E73: out_word = 8'h22;
		16'h1E74: out_word = 8'h42;
		16'h1E75: out_word = 8'h5C;
		16'h1E76: out_word = 8'hFD;
		16'h1E77: out_word = 8'h72;
		16'h1E78: out_word = 8'h0A;
		16'h1E79: out_word = 8'hC9;
		16'h1E7A: out_word = 8'hCD;
		16'h1E7B: out_word = 8'h85;
		16'h1E7C: out_word = 8'h1E;
		16'h1E7D: out_word = 8'hED;
		16'h1E7E: out_word = 8'h79;
		16'h1E7F: out_word = 8'hC9;
		16'h1E80: out_word = 8'hCD;
		16'h1E81: out_word = 8'h85;
		16'h1E82: out_word = 8'h1E;
		16'h1E83: out_word = 8'h02;
		16'h1E84: out_word = 8'hC9;
		16'h1E85: out_word = 8'hCD;
		16'h1E86: out_word = 8'hD5;
		16'h1E87: out_word = 8'h2D;
		16'h1E88: out_word = 8'h38;
		16'h1E89: out_word = 8'h15;
		16'h1E8A: out_word = 8'h28;
		16'h1E8B: out_word = 8'h02;
		16'h1E8C: out_word = 8'hED;
		16'h1E8D: out_word = 8'h44;
		16'h1E8E: out_word = 8'hF5;
		16'h1E8F: out_word = 8'hCD;
		16'h1E90: out_word = 8'h99;
		16'h1E91: out_word = 8'h1E;
		16'h1E92: out_word = 8'hF1;
		16'h1E93: out_word = 8'hC9;
		16'h1E94: out_word = 8'hCD;
		16'h1E95: out_word = 8'hD5;
		16'h1E96: out_word = 8'h2D;
		16'h1E97: out_word = 8'h18;
		16'h1E98: out_word = 8'h03;
		16'h1E99: out_word = 8'hCD;
		16'h1E9A: out_word = 8'hA2;
		16'h1E9B: out_word = 8'h2D;
		16'h1E9C: out_word = 8'h38;
		16'h1E9D: out_word = 8'h01;
		16'h1E9E: out_word = 8'hC8;
		16'h1E9F: out_word = 8'hCF;
		16'h1EA0: out_word = 8'h0A;
		16'h1EA1: out_word = 8'hCD;
		16'h1EA2: out_word = 8'h67;
		16'h1EA3: out_word = 8'h1E;
		16'h1EA4: out_word = 8'h01;
		16'h1EA5: out_word = 8'h00;
		16'h1EA6: out_word = 8'h00;
		16'h1EA7: out_word = 8'hCD;
		16'h1EA8: out_word = 8'h45;
		16'h1EA9: out_word = 8'h1E;
		16'h1EAA: out_word = 8'h18;
		16'h1EAB: out_word = 8'h03;
		16'h1EAC: out_word = 8'hCD;
		16'h1EAD: out_word = 8'h99;
		16'h1EAE: out_word = 8'h1E;
		16'h1EAF: out_word = 8'h78;
		16'h1EB0: out_word = 8'hB1;
		16'h1EB1: out_word = 8'h20;
		16'h1EB2: out_word = 8'h04;
		16'h1EB3: out_word = 8'hED;
		16'h1EB4: out_word = 8'h4B;
		16'h1EB5: out_word = 8'hB2;
		16'h1EB6: out_word = 8'h5C;
		16'h1EB7: out_word = 8'hC5;
		16'h1EB8: out_word = 8'hED;
		16'h1EB9: out_word = 8'h5B;
		16'h1EBA: out_word = 8'h4B;
		16'h1EBB: out_word = 8'h5C;
		16'h1EBC: out_word = 8'h2A;
		16'h1EBD: out_word = 8'h59;
		16'h1EBE: out_word = 8'h5C;
		16'h1EBF: out_word = 8'h2B;
		16'h1EC0: out_word = 8'hCD;
		16'h1EC1: out_word = 8'hE5;
		16'h1EC2: out_word = 8'h19;
		16'h1EC3: out_word = 8'hCD;
		16'h1EC4: out_word = 8'h6B;
		16'h1EC5: out_word = 8'h0D;
		16'h1EC6: out_word = 8'h2A;
		16'h1EC7: out_word = 8'h65;
		16'h1EC8: out_word = 8'h5C;
		16'h1EC9: out_word = 8'h11;
		16'h1ECA: out_word = 8'h32;
		16'h1ECB: out_word = 8'h00;
		16'h1ECC: out_word = 8'h19;
		16'h1ECD: out_word = 8'hD1;
		16'h1ECE: out_word = 8'hED;
		16'h1ECF: out_word = 8'h52;
		16'h1ED0: out_word = 8'h30;
		16'h1ED1: out_word = 8'h08;
		16'h1ED2: out_word = 8'h2A;
		16'h1ED3: out_word = 8'hB4;
		16'h1ED4: out_word = 8'h5C;
		16'h1ED5: out_word = 8'hA7;
		16'h1ED6: out_word = 8'hED;
		16'h1ED7: out_word = 8'h52;
		16'h1ED8: out_word = 8'h30;
		16'h1ED9: out_word = 8'h02;
		16'h1EDA: out_word = 8'hCF;
		16'h1EDB: out_word = 8'h15;
		16'h1EDC: out_word = 8'hEB;
		16'h1EDD: out_word = 8'h22;
		16'h1EDE: out_word = 8'hB2;
		16'h1EDF: out_word = 8'h5C;
		16'h1EE0: out_word = 8'hD1;
		16'h1EE1: out_word = 8'hC1;
		16'h1EE2: out_word = 8'h36;
		16'h1EE3: out_word = 8'h3E;
		16'h1EE4: out_word = 8'h2B;
		16'h1EE5: out_word = 8'hF9;
		16'h1EE6: out_word = 8'hC5;
		16'h1EE7: out_word = 8'hED;
		16'h1EE8: out_word = 8'h73;
		16'h1EE9: out_word = 8'h3D;
		16'h1EEA: out_word = 8'h5C;
		16'h1EEB: out_word = 8'hEB;
		16'h1EEC: out_word = 8'hE9;
		16'h1EED: out_word = 8'hD1;
		16'h1EEE: out_word = 8'hFD;
		16'h1EEF: out_word = 8'h66;
		16'h1EF0: out_word = 8'h0D;
		16'h1EF1: out_word = 8'h24;
		16'h1EF2: out_word = 8'hE3;
		16'h1EF3: out_word = 8'h33;
		16'h1EF4: out_word = 8'hED;
		16'h1EF5: out_word = 8'h4B;
		16'h1EF6: out_word = 8'h45;
		16'h1EF7: out_word = 8'h5C;
		16'h1EF8: out_word = 8'hC5;
		16'h1EF9: out_word = 8'hE5;
		16'h1EFA: out_word = 8'hED;
		16'h1EFB: out_word = 8'h73;
		16'h1EFC: out_word = 8'h3D;
		16'h1EFD: out_word = 8'h5C;
		16'h1EFE: out_word = 8'hD5;
		16'h1EFF: out_word = 8'hCD;
		16'h1F00: out_word = 8'h67;
		16'h1F01: out_word = 8'h1E;
		16'h1F02: out_word = 8'h01;
		16'h1F03: out_word = 8'h14;
		16'h1F04: out_word = 8'h00;
		16'h1F05: out_word = 8'h2A;
		16'h1F06: out_word = 8'h65;
		16'h1F07: out_word = 8'h5C;
		16'h1F08: out_word = 8'h09;
		16'h1F09: out_word = 8'h38;
		16'h1F0A: out_word = 8'h0A;
		16'h1F0B: out_word = 8'hEB;
		16'h1F0C: out_word = 8'h21;
		16'h1F0D: out_word = 8'h50;
		16'h1F0E: out_word = 8'h00;
		16'h1F0F: out_word = 8'h19;
		16'h1F10: out_word = 8'h38;
		16'h1F11: out_word = 8'h03;
		16'h1F12: out_word = 8'hED;
		16'h1F13: out_word = 8'h72;
		16'h1F14: out_word = 8'hD8;
		16'h1F15: out_word = 8'h2E;
		16'h1F16: out_word = 8'h03;
		16'h1F17: out_word = 8'hC3;
		16'h1F18: out_word = 8'h55;
		16'h1F19: out_word = 8'h00;
		16'h1F1A: out_word = 8'h01;
		16'h1F1B: out_word = 8'h00;
		16'h1F1C: out_word = 8'h00;
		16'h1F1D: out_word = 8'hCD;
		16'h1F1E: out_word = 8'h05;
		16'h1F1F: out_word = 8'h1F;
		16'h1F20: out_word = 8'h44;
		16'h1F21: out_word = 8'h4D;
		16'h1F22: out_word = 8'hC9;
		16'h1F23: out_word = 8'hC1;
		16'h1F24: out_word = 8'hE1;
		16'h1F25: out_word = 8'hD1;
		16'h1F26: out_word = 8'h7A;
		16'h1F27: out_word = 8'hFE;
		16'h1F28: out_word = 8'h3E;
		16'h1F29: out_word = 8'h28;
		16'h1F2A: out_word = 8'h0B;
		16'h1F2B: out_word = 8'h3B;
		16'h1F2C: out_word = 8'hE3;
		16'h1F2D: out_word = 8'hEB;
		16'h1F2E: out_word = 8'hED;
		16'h1F2F: out_word = 8'h73;
		16'h1F30: out_word = 8'h3D;
		16'h1F31: out_word = 8'h5C;
		16'h1F32: out_word = 8'hC5;
		16'h1F33: out_word = 8'hC3;
		16'h1F34: out_word = 8'h73;
		16'h1F35: out_word = 8'h1E;
		16'h1F36: out_word = 8'hD5;
		16'h1F37: out_word = 8'hE5;
		16'h1F38: out_word = 8'hCF;
		16'h1F39: out_word = 8'h06;
		16'h1F3A: out_word = 8'hCD;
		16'h1F3B: out_word = 8'h99;
		16'h1F3C: out_word = 8'h1E;
		16'h1F3D: out_word = 8'h76;
		16'h1F3E: out_word = 8'h0B;
		16'h1F3F: out_word = 8'h78;
		16'h1F40: out_word = 8'hB1;
		16'h1F41: out_word = 8'h28;
		16'h1F42: out_word = 8'h0C;
		16'h1F43: out_word = 8'h78;
		16'h1F44: out_word = 8'hA1;
		16'h1F45: out_word = 8'h3C;
		16'h1F46: out_word = 8'h20;
		16'h1F47: out_word = 8'h01;
		16'h1F48: out_word = 8'h03;
		16'h1F49: out_word = 8'hFD;
		16'h1F4A: out_word = 8'hCB;
		16'h1F4B: out_word = 8'h01;
		16'h1F4C: out_word = 8'h6E;
		16'h1F4D: out_word = 8'h28;
		16'h1F4E: out_word = 8'hEE;
		16'h1F4F: out_word = 8'hFD;
		16'h1F50: out_word = 8'hCB;
		16'h1F51: out_word = 8'h01;
		16'h1F52: out_word = 8'hAE;
		16'h1F53: out_word = 8'hC9;
		16'h1F54: out_word = 8'h3E;
		16'h1F55: out_word = 8'h7F;
		16'h1F56: out_word = 8'hDB;
		16'h1F57: out_word = 8'hFE;
		16'h1F58: out_word = 8'h1F;
		16'h1F59: out_word = 8'hD8;
		16'h1F5A: out_word = 8'h3E;
		16'h1F5B: out_word = 8'hFE;
		16'h1F5C: out_word = 8'hDB;
		16'h1F5D: out_word = 8'hFE;
		16'h1F5E: out_word = 8'h1F;
		16'h1F5F: out_word = 8'hC9;
		16'h1F60: out_word = 8'hCD;
		16'h1F61: out_word = 8'h30;
		16'h1F62: out_word = 8'h25;
		16'h1F63: out_word = 8'h28;
		16'h1F64: out_word = 8'h05;
		16'h1F65: out_word = 8'h3E;
		16'h1F66: out_word = 8'hCE;
		16'h1F67: out_word = 8'hC3;
		16'h1F68: out_word = 8'h39;
		16'h1F69: out_word = 8'h1E;
		16'h1F6A: out_word = 8'hFD;
		16'h1F6B: out_word = 8'hCB;
		16'h1F6C: out_word = 8'h01;
		16'h1F6D: out_word = 8'hF6;
		16'h1F6E: out_word = 8'hCD;
		16'h1F6F: out_word = 8'h8D;
		16'h1F70: out_word = 8'h2C;
		16'h1F71: out_word = 8'h30;
		16'h1F72: out_word = 8'h16;
		16'h1F73: out_word = 8'hE7;
		16'h1F74: out_word = 8'hFE;
		16'h1F75: out_word = 8'h24;
		16'h1F76: out_word = 8'h20;
		16'h1F77: out_word = 8'h05;
		16'h1F78: out_word = 8'hFD;
		16'h1F79: out_word = 8'hCB;
		16'h1F7A: out_word = 8'h01;
		16'h1F7B: out_word = 8'hB6;
		16'h1F7C: out_word = 8'hE7;
		16'h1F7D: out_word = 8'hFE;
		16'h1F7E: out_word = 8'h28;
		16'h1F7F: out_word = 8'h20;
		16'h1F80: out_word = 8'h3C;
		16'h1F81: out_word = 8'hE7;
		16'h1F82: out_word = 8'hFE;
		16'h1F83: out_word = 8'h29;
		16'h1F84: out_word = 8'h28;
		16'h1F85: out_word = 8'h20;
		16'h1F86: out_word = 8'hCD;
		16'h1F87: out_word = 8'h8D;
		16'h1F88: out_word = 8'h2C;
		16'h1F89: out_word = 8'hD2;
		16'h1F8A: out_word = 8'h8A;
		16'h1F8B: out_word = 8'h1C;
		16'h1F8C: out_word = 8'hEB;
		16'h1F8D: out_word = 8'hE7;
		16'h1F8E: out_word = 8'hFE;
		16'h1F8F: out_word = 8'h24;
		16'h1F90: out_word = 8'h20;
		16'h1F91: out_word = 8'h02;
		16'h1F92: out_word = 8'hEB;
		16'h1F93: out_word = 8'hE7;
		16'h1F94: out_word = 8'hEB;
		16'h1F95: out_word = 8'h01;
		16'h1F96: out_word = 8'h06;
		16'h1F97: out_word = 8'h00;
		16'h1F98: out_word = 8'hCD;
		16'h1F99: out_word = 8'h55;
		16'h1F9A: out_word = 8'h16;
		16'h1F9B: out_word = 8'h23;
		16'h1F9C: out_word = 8'h23;
		16'h1F9D: out_word = 8'h36;
		16'h1F9E: out_word = 8'h0E;
		16'h1F9F: out_word = 8'hFE;
		16'h1FA0: out_word = 8'h2C;
		16'h1FA1: out_word = 8'h20;
		16'h1FA2: out_word = 8'h03;
		16'h1FA3: out_word = 8'hE7;
		16'h1FA4: out_word = 8'h18;
		16'h1FA5: out_word = 8'hE0;
		16'h1FA6: out_word = 8'hFE;
		16'h1FA7: out_word = 8'h29;
		16'h1FA8: out_word = 8'h20;
		16'h1FA9: out_word = 8'h13;
		16'h1FAA: out_word = 8'hE7;
		16'h1FAB: out_word = 8'hFE;
		16'h1FAC: out_word = 8'h3D;
		16'h1FAD: out_word = 8'h20;
		16'h1FAE: out_word = 8'h0E;
		16'h1FAF: out_word = 8'hE7;
		16'h1FB0: out_word = 8'h3A;
		16'h1FB1: out_word = 8'h3B;
		16'h1FB2: out_word = 8'h5C;
		16'h1FB3: out_word = 8'hF5;
		16'h1FB4: out_word = 8'hCD;
		16'h1FB5: out_word = 8'hFB;
		16'h1FB6: out_word = 8'h24;
		16'h1FB7: out_word = 8'hF1;
		16'h1FB8: out_word = 8'hFD;
		16'h1FB9: out_word = 8'hAE;
		16'h1FBA: out_word = 8'h01;
		16'h1FBB: out_word = 8'hE6;
		16'h1FBC: out_word = 8'h40;
		16'h1FBD: out_word = 8'hC2;
		16'h1FBE: out_word = 8'h8A;
		16'h1FBF: out_word = 8'h1C;
		16'h1FC0: out_word = 8'hCD;
		16'h1FC1: out_word = 8'hEE;
		16'h1FC2: out_word = 8'h1B;
		16'h1FC3: out_word = 8'hCD;
		16'h1FC4: out_word = 8'h30;
		16'h1FC5: out_word = 8'h25;
		16'h1FC6: out_word = 8'hE1;
		16'h1FC7: out_word = 8'hC8;
		16'h1FC8: out_word = 8'hE9;
		16'h1FC9: out_word = 8'h3E;
		16'h1FCA: out_word = 8'h03;
		16'h1FCB: out_word = 8'h18;
		16'h1FCC: out_word = 8'h02;
		16'h1FCD: out_word = 8'h3E;
		16'h1FCE: out_word = 8'h02;
		16'h1FCF: out_word = 8'hCD;
		16'h1FD0: out_word = 8'h30;
		16'h1FD1: out_word = 8'h25;
		16'h1FD2: out_word = 8'hC4;
		16'h1FD3: out_word = 8'h01;
		16'h1FD4: out_word = 8'h16;
		16'h1FD5: out_word = 8'hCD;
		16'h1FD6: out_word = 8'h4D;
		16'h1FD7: out_word = 8'h0D;
		16'h1FD8: out_word = 8'hCD;
		16'h1FD9: out_word = 8'hDF;
		16'h1FDA: out_word = 8'h1F;
		16'h1FDB: out_word = 8'hCD;
		16'h1FDC: out_word = 8'hEE;
		16'h1FDD: out_word = 8'h1B;
		16'h1FDE: out_word = 8'hC9;
		16'h1FDF: out_word = 8'hDF;
		16'h1FE0: out_word = 8'hCD;
		16'h1FE1: out_word = 8'h45;
		16'h1FE2: out_word = 8'h20;
		16'h1FE3: out_word = 8'h28;
		16'h1FE4: out_word = 8'h0D;
		16'h1FE5: out_word = 8'hCD;
		16'h1FE6: out_word = 8'h4E;
		16'h1FE7: out_word = 8'h20;
		16'h1FE8: out_word = 8'h28;
		16'h1FE9: out_word = 8'hFB;
		16'h1FEA: out_word = 8'hCD;
		16'h1FEB: out_word = 8'hFC;
		16'h1FEC: out_word = 8'h1F;
		16'h1FED: out_word = 8'hCD;
		16'h1FEE: out_word = 8'h4E;
		16'h1FEF: out_word = 8'h20;
		16'h1FF0: out_word = 8'h28;
		16'h1FF1: out_word = 8'hF3;
		16'h1FF2: out_word = 8'hFE;
		16'h1FF3: out_word = 8'h29;
		16'h1FF4: out_word = 8'hC8;
		16'h1FF5: out_word = 8'hCD;
		16'h1FF6: out_word = 8'hC3;
		16'h1FF7: out_word = 8'h1F;
		16'h1FF8: out_word = 8'h3E;
		16'h1FF9: out_word = 8'h0D;
		16'h1FFA: out_word = 8'hD7;
		16'h1FFB: out_word = 8'hC9;
		16'h1FFC: out_word = 8'hDF;
		16'h1FFD: out_word = 8'hFE;
		16'h1FFE: out_word = 8'hAC;
		16'h1FFF: out_word = 8'h20;
		16'h2000: out_word = 8'h0D;
		16'h2001: out_word = 8'hCD;
		16'h2002: out_word = 8'h79;
		16'h2003: out_word = 8'h1C;
		16'h2004: out_word = 8'hCD;
		16'h2005: out_word = 8'hC3;
		16'h2006: out_word = 8'h1F;
		16'h2007: out_word = 8'hCD;
		16'h2008: out_word = 8'h07;
		16'h2009: out_word = 8'h23;
		16'h200A: out_word = 8'h3E;
		16'h200B: out_word = 8'h16;
		16'h200C: out_word = 8'h18;
		16'h200D: out_word = 8'h10;
		16'h200E: out_word = 8'hFE;
		16'h200F: out_word = 8'hAD;
		16'h2010: out_word = 8'h20;
		16'h2011: out_word = 8'h12;
		16'h2012: out_word = 8'hE7;
		16'h2013: out_word = 8'hCD;
		16'h2014: out_word = 8'h82;
		16'h2015: out_word = 8'h1C;
		16'h2016: out_word = 8'hCD;
		16'h2017: out_word = 8'hC3;
		16'h2018: out_word = 8'h1F;
		16'h2019: out_word = 8'hCD;
		16'h201A: out_word = 8'h99;
		16'h201B: out_word = 8'h1E;
		16'h201C: out_word = 8'h3E;
		16'h201D: out_word = 8'h17;
		16'h201E: out_word = 8'hD7;
		16'h201F: out_word = 8'h79;
		16'h2020: out_word = 8'hD7;
		16'h2021: out_word = 8'h78;
		16'h2022: out_word = 8'hD7;
		16'h2023: out_word = 8'hC9;
		16'h2024: out_word = 8'hCD;
		16'h2025: out_word = 8'hF2;
		16'h2026: out_word = 8'h21;
		16'h2027: out_word = 8'hD0;
		16'h2028: out_word = 8'hCD;
		16'h2029: out_word = 8'h70;
		16'h202A: out_word = 8'h20;
		16'h202B: out_word = 8'hD0;
		16'h202C: out_word = 8'hCD;
		16'h202D: out_word = 8'hFB;
		16'h202E: out_word = 8'h24;
		16'h202F: out_word = 8'hCD;
		16'h2030: out_word = 8'hC3;
		16'h2031: out_word = 8'h1F;
		16'h2032: out_word = 8'hFD;
		16'h2033: out_word = 8'hCB;
		16'h2034: out_word = 8'h01;
		16'h2035: out_word = 8'h76;
		16'h2036: out_word = 8'hCC;
		16'h2037: out_word = 8'hF1;
		16'h2038: out_word = 8'h2B;
		16'h2039: out_word = 8'hC2;
		16'h203A: out_word = 8'hE3;
		16'h203B: out_word = 8'h2D;
		16'h203C: out_word = 8'h78;
		16'h203D: out_word = 8'hB1;
		16'h203E: out_word = 8'h0B;
		16'h203F: out_word = 8'hC8;
		16'h2040: out_word = 8'h1A;
		16'h2041: out_word = 8'h13;
		16'h2042: out_word = 8'hD7;
		16'h2043: out_word = 8'h18;
		16'h2044: out_word = 8'hF7;
		16'h2045: out_word = 8'hFE;
		16'h2046: out_word = 8'h29;
		16'h2047: out_word = 8'hC8;
		16'h2048: out_word = 8'hFE;
		16'h2049: out_word = 8'h0D;
		16'h204A: out_word = 8'hC8;
		16'h204B: out_word = 8'hFE;
		16'h204C: out_word = 8'h3A;
		16'h204D: out_word = 8'hC9;
		16'h204E: out_word = 8'hDF;
		16'h204F: out_word = 8'hFE;
		16'h2050: out_word = 8'h3B;
		16'h2051: out_word = 8'h28;
		16'h2052: out_word = 8'h14;
		16'h2053: out_word = 8'hFE;
		16'h2054: out_word = 8'h2C;
		16'h2055: out_word = 8'h20;
		16'h2056: out_word = 8'h0A;
		16'h2057: out_word = 8'hCD;
		16'h2058: out_word = 8'h30;
		16'h2059: out_word = 8'h25;
		16'h205A: out_word = 8'h28;
		16'h205B: out_word = 8'h0B;
		16'h205C: out_word = 8'h3E;
		16'h205D: out_word = 8'h06;
		16'h205E: out_word = 8'hD7;
		16'h205F: out_word = 8'h18;
		16'h2060: out_word = 8'h06;
		16'h2061: out_word = 8'hFE;
		16'h2062: out_word = 8'h27;
		16'h2063: out_word = 8'hC0;
		16'h2064: out_word = 8'hCD;
		16'h2065: out_word = 8'hF5;
		16'h2066: out_word = 8'h1F;
		16'h2067: out_word = 8'hE7;
		16'h2068: out_word = 8'hCD;
		16'h2069: out_word = 8'h45;
		16'h206A: out_word = 8'h20;
		16'h206B: out_word = 8'h20;
		16'h206C: out_word = 8'h01;
		16'h206D: out_word = 8'hC1;
		16'h206E: out_word = 8'hBF;
		16'h206F: out_word = 8'hC9;
		16'h2070: out_word = 8'hFE;
		16'h2071: out_word = 8'h23;
		16'h2072: out_word = 8'h37;
		16'h2073: out_word = 8'hC0;
		16'h2074: out_word = 8'hE7;
		16'h2075: out_word = 8'hCD;
		16'h2076: out_word = 8'h82;
		16'h2077: out_word = 8'h1C;
		16'h2078: out_word = 8'hA7;
		16'h2079: out_word = 8'hCD;
		16'h207A: out_word = 8'hC3;
		16'h207B: out_word = 8'h1F;
		16'h207C: out_word = 8'hCD;
		16'h207D: out_word = 8'h94;
		16'h207E: out_word = 8'h1E;
		16'h207F: out_word = 8'hFE;
		16'h2080: out_word = 8'h10;
		16'h2081: out_word = 8'hD2;
		16'h2082: out_word = 8'h0E;
		16'h2083: out_word = 8'h16;
		16'h2084: out_word = 8'hCD;
		16'h2085: out_word = 8'h01;
		16'h2086: out_word = 8'h16;
		16'h2087: out_word = 8'hA7;
		16'h2088: out_word = 8'hC9;
		16'h2089: out_word = 8'hCD;
		16'h208A: out_word = 8'h30;
		16'h208B: out_word = 8'h25;
		16'h208C: out_word = 8'h28;
		16'h208D: out_word = 8'h08;
		16'h208E: out_word = 8'h3E;
		16'h208F: out_word = 8'h01;
		16'h2090: out_word = 8'hCD;
		16'h2091: out_word = 8'h01;
		16'h2092: out_word = 8'h16;
		16'h2093: out_word = 8'hCD;
		16'h2094: out_word = 8'h6E;
		16'h2095: out_word = 8'h0D;
		16'h2096: out_word = 8'hFD;
		16'h2097: out_word = 8'h36;
		16'h2098: out_word = 8'h02;
		16'h2099: out_word = 8'h01;
		16'h209A: out_word = 8'hCD;
		16'h209B: out_word = 8'hC1;
		16'h209C: out_word = 8'h20;
		16'h209D: out_word = 8'hCD;
		16'h209E: out_word = 8'hEE;
		16'h209F: out_word = 8'h1B;
		16'h20A0: out_word = 8'hED;
		16'h20A1: out_word = 8'h4B;
		16'h20A2: out_word = 8'h88;
		16'h20A3: out_word = 8'h5C;
		16'h20A4: out_word = 8'h3A;
		16'h20A5: out_word = 8'h6B;
		16'h20A6: out_word = 8'h5C;
		16'h20A7: out_word = 8'hB8;
		16'h20A8: out_word = 8'h38;
		16'h20A9: out_word = 8'h03;
		16'h20AA: out_word = 8'h0E;
		16'h20AB: out_word = 8'h21;
		16'h20AC: out_word = 8'h47;
		16'h20AD: out_word = 8'hED;
		16'h20AE: out_word = 8'h43;
		16'h20AF: out_word = 8'h88;
		16'h20B0: out_word = 8'h5C;
		16'h20B1: out_word = 8'h3E;
		16'h20B2: out_word = 8'h19;
		16'h20B3: out_word = 8'h90;
		16'h20B4: out_word = 8'h32;
		16'h20B5: out_word = 8'h8C;
		16'h20B6: out_word = 8'h5C;
		16'h20B7: out_word = 8'hFD;
		16'h20B8: out_word = 8'hCB;
		16'h20B9: out_word = 8'h02;
		16'h20BA: out_word = 8'h86;
		16'h20BB: out_word = 8'hCD;
		16'h20BC: out_word = 8'hD9;
		16'h20BD: out_word = 8'h0D;
		16'h20BE: out_word = 8'hC3;
		16'h20BF: out_word = 8'h6E;
		16'h20C0: out_word = 8'h0D;
		16'h20C1: out_word = 8'hCD;
		16'h20C2: out_word = 8'h4E;
		16'h20C3: out_word = 8'h20;
		16'h20C4: out_word = 8'h28;
		16'h20C5: out_word = 8'hFB;
		16'h20C6: out_word = 8'hFE;
		16'h20C7: out_word = 8'h28;
		16'h20C8: out_word = 8'h20;
		16'h20C9: out_word = 8'h0E;
		16'h20CA: out_word = 8'hE7;
		16'h20CB: out_word = 8'hCD;
		16'h20CC: out_word = 8'hDF;
		16'h20CD: out_word = 8'h1F;
		16'h20CE: out_word = 8'hDF;
		16'h20CF: out_word = 8'hFE;
		16'h20D0: out_word = 8'h29;
		16'h20D1: out_word = 8'hC2;
		16'h20D2: out_word = 8'h8A;
		16'h20D3: out_word = 8'h1C;
		16'h20D4: out_word = 8'hE7;
		16'h20D5: out_word = 8'hC3;
		16'h20D6: out_word = 8'hB2;
		16'h20D7: out_word = 8'h21;
		16'h20D8: out_word = 8'hFE;
		16'h20D9: out_word = 8'hCA;
		16'h20DA: out_word = 8'h20;
		16'h20DB: out_word = 8'h11;
		16'h20DC: out_word = 8'hE7;
		16'h20DD: out_word = 8'hCD;
		16'h20DE: out_word = 8'h1F;
		16'h20DF: out_word = 8'h1C;
		16'h20E0: out_word = 8'hFD;
		16'h20E1: out_word = 8'hCB;
		16'h20E2: out_word = 8'h37;
		16'h20E3: out_word = 8'hFE;
		16'h20E4: out_word = 8'hFD;
		16'h20E5: out_word = 8'hCB;
		16'h20E6: out_word = 8'h01;
		16'h20E7: out_word = 8'h76;
		16'h20E8: out_word = 8'hC2;
		16'h20E9: out_word = 8'h8A;
		16'h20EA: out_word = 8'h1C;
		16'h20EB: out_word = 8'h18;
		16'h20EC: out_word = 8'h0D;
		16'h20ED: out_word = 8'hCD;
		16'h20EE: out_word = 8'h8D;
		16'h20EF: out_word = 8'h2C;
		16'h20F0: out_word = 8'hD2;
		16'h20F1: out_word = 8'hAF;
		16'h20F2: out_word = 8'h21;
		16'h20F3: out_word = 8'hCD;
		16'h20F4: out_word = 8'h1F;
		16'h20F5: out_word = 8'h1C;
		16'h20F6: out_word = 8'hFD;
		16'h20F7: out_word = 8'hCB;
		16'h20F8: out_word = 8'h37;
		16'h20F9: out_word = 8'hBE;
		16'h20FA: out_word = 8'hCD;
		16'h20FB: out_word = 8'h30;
		16'h20FC: out_word = 8'h25;
		16'h20FD: out_word = 8'hCA;
		16'h20FE: out_word = 8'hB2;
		16'h20FF: out_word = 8'h21;
		16'h2100: out_word = 8'hCD;
		16'h2101: out_word = 8'hBF;
		16'h2102: out_word = 8'h16;
		16'h2103: out_word = 8'h21;
		16'h2104: out_word = 8'h71;
		16'h2105: out_word = 8'h5C;
		16'h2106: out_word = 8'hCB;
		16'h2107: out_word = 8'hB6;
		16'h2108: out_word = 8'hCB;
		16'h2109: out_word = 8'hEE;
		16'h210A: out_word = 8'h01;
		16'h210B: out_word = 8'h01;
		16'h210C: out_word = 8'h00;
		16'h210D: out_word = 8'hCB;
		16'h210E: out_word = 8'h7E;
		16'h210F: out_word = 8'h20;
		16'h2110: out_word = 8'h0B;
		16'h2111: out_word = 8'h3A;
		16'h2112: out_word = 8'h3B;
		16'h2113: out_word = 8'h5C;
		16'h2114: out_word = 8'hE6;
		16'h2115: out_word = 8'h40;
		16'h2116: out_word = 8'h20;
		16'h2117: out_word = 8'h02;
		16'h2118: out_word = 8'h0E;
		16'h2119: out_word = 8'h03;
		16'h211A: out_word = 8'hB6;
		16'h211B: out_word = 8'h77;
		16'h211C: out_word = 8'hF7;
		16'h211D: out_word = 8'h36;
		16'h211E: out_word = 8'h0D;
		16'h211F: out_word = 8'h79;
		16'h2120: out_word = 8'h0F;
		16'h2121: out_word = 8'h0F;
		16'h2122: out_word = 8'h30;
		16'h2123: out_word = 8'h05;
		16'h2124: out_word = 8'h3E;
		16'h2125: out_word = 8'h22;
		16'h2126: out_word = 8'h12;
		16'h2127: out_word = 8'h2B;
		16'h2128: out_word = 8'h77;
		16'h2129: out_word = 8'h22;
		16'h212A: out_word = 8'h5B;
		16'h212B: out_word = 8'h5C;
		16'h212C: out_word = 8'hFD;
		16'h212D: out_word = 8'hCB;
		16'h212E: out_word = 8'h37;
		16'h212F: out_word = 8'h7E;
		16'h2130: out_word = 8'h20;
		16'h2131: out_word = 8'h2C;
		16'h2132: out_word = 8'h2A;
		16'h2133: out_word = 8'h5D;
		16'h2134: out_word = 8'h5C;
		16'h2135: out_word = 8'hE5;
		16'h2136: out_word = 8'h2A;
		16'h2137: out_word = 8'h3D;
		16'h2138: out_word = 8'h5C;
		16'h2139: out_word = 8'hE5;
		16'h213A: out_word = 8'h21;
		16'h213B: out_word = 8'h3A;
		16'h213C: out_word = 8'h21;
		16'h213D: out_word = 8'hE5;
		16'h213E: out_word = 8'hFD;
		16'h213F: out_word = 8'hCB;
		16'h2140: out_word = 8'h30;
		16'h2141: out_word = 8'h66;
		16'h2142: out_word = 8'h28;
		16'h2143: out_word = 8'h04;
		16'h2144: out_word = 8'hED;
		16'h2145: out_word = 8'h73;
		16'h2146: out_word = 8'h3D;
		16'h2147: out_word = 8'h5C;
		16'h2148: out_word = 8'h2A;
		16'h2149: out_word = 8'h61;
		16'h214A: out_word = 8'h5C;
		16'h214B: out_word = 8'hCD;
		16'h214C: out_word = 8'hA7;
		16'h214D: out_word = 8'h11;
		16'h214E: out_word = 8'hFD;
		16'h214F: out_word = 8'h36;
		16'h2150: out_word = 8'h00;
		16'h2151: out_word = 8'hFF;
		16'h2152: out_word = 8'hCD;
		16'h2153: out_word = 8'h2C;
		16'h2154: out_word = 8'h0F;
		16'h2155: out_word = 8'hFD;
		16'h2156: out_word = 8'hCB;
		16'h2157: out_word = 8'h01;
		16'h2158: out_word = 8'hBE;
		16'h2159: out_word = 8'hCD;
		16'h215A: out_word = 8'hB9;
		16'h215B: out_word = 8'h21;
		16'h215C: out_word = 8'h18;
		16'h215D: out_word = 8'h03;
		16'h215E: out_word = 8'hCD;
		16'h215F: out_word = 8'h2C;
		16'h2160: out_word = 8'h0F;
		16'h2161: out_word = 8'hFD;
		16'h2162: out_word = 8'h36;
		16'h2163: out_word = 8'h22;
		16'h2164: out_word = 8'h00;
		16'h2165: out_word = 8'hCD;
		16'h2166: out_word = 8'hD6;
		16'h2167: out_word = 8'h21;
		16'h2168: out_word = 8'h20;
		16'h2169: out_word = 8'h0A;
		16'h216A: out_word = 8'hCD;
		16'h216B: out_word = 8'h1D;
		16'h216C: out_word = 8'h11;
		16'h216D: out_word = 8'hED;
		16'h216E: out_word = 8'h4B;
		16'h216F: out_word = 8'h82;
		16'h2170: out_word = 8'h5C;
		16'h2171: out_word = 8'hCD;
		16'h2172: out_word = 8'hD9;
		16'h2173: out_word = 8'h0D;
		16'h2174: out_word = 8'h21;
		16'h2175: out_word = 8'h71;
		16'h2176: out_word = 8'h5C;
		16'h2177: out_word = 8'hCB;
		16'h2178: out_word = 8'hAE;
		16'h2179: out_word = 8'hCB;
		16'h217A: out_word = 8'h7E;
		16'h217B: out_word = 8'hCB;
		16'h217C: out_word = 8'hBE;
		16'h217D: out_word = 8'h20;
		16'h217E: out_word = 8'h1C;
		16'h217F: out_word = 8'hE1;
		16'h2180: out_word = 8'hE1;
		16'h2181: out_word = 8'h22;
		16'h2182: out_word = 8'h3D;
		16'h2183: out_word = 8'h5C;
		16'h2184: out_word = 8'hE1;
		16'h2185: out_word = 8'h22;
		16'h2186: out_word = 8'h5F;
		16'h2187: out_word = 8'h5C;
		16'h2188: out_word = 8'hFD;
		16'h2189: out_word = 8'hCB;
		16'h218A: out_word = 8'h01;
		16'h218B: out_word = 8'hFE;
		16'h218C: out_word = 8'hCD;
		16'h218D: out_word = 8'hB9;
		16'h218E: out_word = 8'h21;
		16'h218F: out_word = 8'h2A;
		16'h2190: out_word = 8'h5F;
		16'h2191: out_word = 8'h5C;
		16'h2192: out_word = 8'hFD;
		16'h2193: out_word = 8'h36;
		16'h2194: out_word = 8'h26;
		16'h2195: out_word = 8'h00;
		16'h2196: out_word = 8'h22;
		16'h2197: out_word = 8'h5D;
		16'h2198: out_word = 8'h5C;
		16'h2199: out_word = 8'h18;
		16'h219A: out_word = 8'h17;
		16'h219B: out_word = 8'h2A;
		16'h219C: out_word = 8'h63;
		16'h219D: out_word = 8'h5C;
		16'h219E: out_word = 8'hED;
		16'h219F: out_word = 8'h5B;
		16'h21A0: out_word = 8'h61;
		16'h21A1: out_word = 8'h5C;
		16'h21A2: out_word = 8'h37;
		16'h21A3: out_word = 8'hED;
		16'h21A4: out_word = 8'h52;
		16'h21A5: out_word = 8'h44;
		16'h21A6: out_word = 8'h4D;
		16'h21A7: out_word = 8'hCD;
		16'h21A8: out_word = 8'hB2;
		16'h21A9: out_word = 8'h2A;
		16'h21AA: out_word = 8'hCD;
		16'h21AB: out_word = 8'hFF;
		16'h21AC: out_word = 8'h2A;
		16'h21AD: out_word = 8'h18;
		16'h21AE: out_word = 8'h03;
		16'h21AF: out_word = 8'hCD;
		16'h21B0: out_word = 8'hFC;
		16'h21B1: out_word = 8'h1F;
		16'h21B2: out_word = 8'hCD;
		16'h21B3: out_word = 8'h4E;
		16'h21B4: out_word = 8'h20;
		16'h21B5: out_word = 8'hCA;
		16'h21B6: out_word = 8'hC1;
		16'h21B7: out_word = 8'h20;
		16'h21B8: out_word = 8'hC9;
		16'h21B9: out_word = 8'h2A;
		16'h21BA: out_word = 8'h61;
		16'h21BB: out_word = 8'h5C;
		16'h21BC: out_word = 8'h22;
		16'h21BD: out_word = 8'h5D;
		16'h21BE: out_word = 8'h5C;
		16'h21BF: out_word = 8'hDF;
		16'h21C0: out_word = 8'hFE;
		16'h21C1: out_word = 8'hE2;
		16'h21C2: out_word = 8'h28;
		16'h21C3: out_word = 8'h0C;
		16'h21C4: out_word = 8'h3A;
		16'h21C5: out_word = 8'h71;
		16'h21C6: out_word = 8'h5C;
		16'h21C7: out_word = 8'hCD;
		16'h21C8: out_word = 8'h59;
		16'h21C9: out_word = 8'h1C;
		16'h21CA: out_word = 8'hDF;
		16'h21CB: out_word = 8'hFE;
		16'h21CC: out_word = 8'h0D;
		16'h21CD: out_word = 8'hC8;
		16'h21CE: out_word = 8'hCF;
		16'h21CF: out_word = 8'h0B;
		16'h21D0: out_word = 8'hCD;
		16'h21D1: out_word = 8'h30;
		16'h21D2: out_word = 8'h25;
		16'h21D3: out_word = 8'hC8;
		16'h21D4: out_word = 8'hCF;
		16'h21D5: out_word = 8'h10;
		16'h21D6: out_word = 8'h2A;
		16'h21D7: out_word = 8'h51;
		16'h21D8: out_word = 8'h5C;
		16'h21D9: out_word = 8'h23;
		16'h21DA: out_word = 8'h23;
		16'h21DB: out_word = 8'h23;
		16'h21DC: out_word = 8'h23;
		16'h21DD: out_word = 8'h7E;
		16'h21DE: out_word = 8'hFE;
		16'h21DF: out_word = 8'h4B;
		16'h21E0: out_word = 8'hC9;
		16'h21E1: out_word = 8'hE7;
		16'h21E2: out_word = 8'hCD;
		16'h21E3: out_word = 8'hF2;
		16'h21E4: out_word = 8'h21;
		16'h21E5: out_word = 8'hD8;
		16'h21E6: out_word = 8'hDF;
		16'h21E7: out_word = 8'hFE;
		16'h21E8: out_word = 8'h2C;
		16'h21E9: out_word = 8'h28;
		16'h21EA: out_word = 8'hF6;
		16'h21EB: out_word = 8'hFE;
		16'h21EC: out_word = 8'h3B;
		16'h21ED: out_word = 8'h28;
		16'h21EE: out_word = 8'hF2;
		16'h21EF: out_word = 8'hC3;
		16'h21F0: out_word = 8'h8A;
		16'h21F1: out_word = 8'h1C;
		16'h21F2: out_word = 8'hFE;
		16'h21F3: out_word = 8'hD9;
		16'h21F4: out_word = 8'hD8;
		16'h21F5: out_word = 8'hFE;
		16'h21F6: out_word = 8'hDF;
		16'h21F7: out_word = 8'h3F;
		16'h21F8: out_word = 8'hD8;
		16'h21F9: out_word = 8'hF5;
		16'h21FA: out_word = 8'hE7;
		16'h21FB: out_word = 8'hF1;
		16'h21FC: out_word = 8'hD6;
		16'h21FD: out_word = 8'hC9;
		16'h21FE: out_word = 8'hF5;
		16'h21FF: out_word = 8'hCD;
		16'h2200: out_word = 8'h82;
		16'h2201: out_word = 8'h1C;
		16'h2202: out_word = 8'hF1;
		16'h2203: out_word = 8'hA7;
		16'h2204: out_word = 8'hCD;
		16'h2205: out_word = 8'hC3;
		16'h2206: out_word = 8'h1F;
		16'h2207: out_word = 8'hF5;
		16'h2208: out_word = 8'hCD;
		16'h2209: out_word = 8'h94;
		16'h220A: out_word = 8'h1E;
		16'h220B: out_word = 8'h57;
		16'h220C: out_word = 8'hF1;
		16'h220D: out_word = 8'hD7;
		16'h220E: out_word = 8'h7A;
		16'h220F: out_word = 8'hD7;
		16'h2210: out_word = 8'hC9;
		16'h2211: out_word = 8'hD6;
		16'h2212: out_word = 8'h11;
		16'h2213: out_word = 8'hCE;
		16'h2214: out_word = 8'h00;
		16'h2215: out_word = 8'h28;
		16'h2216: out_word = 8'h1D;
		16'h2217: out_word = 8'hD6;
		16'h2218: out_word = 8'h02;
		16'h2219: out_word = 8'hCE;
		16'h221A: out_word = 8'h00;
		16'h221B: out_word = 8'h28;
		16'h221C: out_word = 8'h56;
		16'h221D: out_word = 8'hFE;
		16'h221E: out_word = 8'h01;
		16'h221F: out_word = 8'h7A;
		16'h2220: out_word = 8'h06;
		16'h2221: out_word = 8'h01;
		16'h2222: out_word = 8'h20;
		16'h2223: out_word = 8'h04;
		16'h2224: out_word = 8'h07;
		16'h2225: out_word = 8'h07;
		16'h2226: out_word = 8'h06;
		16'h2227: out_word = 8'h04;
		16'h2228: out_word = 8'h4F;
		16'h2229: out_word = 8'h7A;
		16'h222A: out_word = 8'hFE;
		16'h222B: out_word = 8'h02;
		16'h222C: out_word = 8'h30;
		16'h222D: out_word = 8'h16;
		16'h222E: out_word = 8'h79;
		16'h222F: out_word = 8'h21;
		16'h2230: out_word = 8'h91;
		16'h2231: out_word = 8'h5C;
		16'h2232: out_word = 8'h18;
		16'h2233: out_word = 8'h38;
		16'h2234: out_word = 8'h7A;
		16'h2235: out_word = 8'h06;
		16'h2236: out_word = 8'h07;
		16'h2237: out_word = 8'h38;
		16'h2238: out_word = 8'h05;
		16'h2239: out_word = 8'h07;
		16'h223A: out_word = 8'h07;
		16'h223B: out_word = 8'h07;
		16'h223C: out_word = 8'h06;
		16'h223D: out_word = 8'h38;
		16'h223E: out_word = 8'h4F;
		16'h223F: out_word = 8'h7A;
		16'h2240: out_word = 8'hFE;
		16'h2241: out_word = 8'h0A;
		16'h2242: out_word = 8'h38;
		16'h2243: out_word = 8'h02;
		16'h2244: out_word = 8'hCF;
		16'h2245: out_word = 8'h13;
		16'h2246: out_word = 8'h21;
		16'h2247: out_word = 8'h8F;
		16'h2248: out_word = 8'h5C;
		16'h2249: out_word = 8'hFE;
		16'h224A: out_word = 8'h08;
		16'h224B: out_word = 8'h38;
		16'h224C: out_word = 8'h0B;
		16'h224D: out_word = 8'h7E;
		16'h224E: out_word = 8'h28;
		16'h224F: out_word = 8'h07;
		16'h2250: out_word = 8'hB0;
		16'h2251: out_word = 8'h2F;
		16'h2252: out_word = 8'hE6;
		16'h2253: out_word = 8'h24;
		16'h2254: out_word = 8'h28;
		16'h2255: out_word = 8'h01;
		16'h2256: out_word = 8'h78;
		16'h2257: out_word = 8'h4F;
		16'h2258: out_word = 8'h79;
		16'h2259: out_word = 8'hCD;
		16'h225A: out_word = 8'h6C;
		16'h225B: out_word = 8'h22;
		16'h225C: out_word = 8'h3E;
		16'h225D: out_word = 8'h07;
		16'h225E: out_word = 8'hBA;
		16'h225F: out_word = 8'h9F;
		16'h2260: out_word = 8'hCD;
		16'h2261: out_word = 8'h6C;
		16'h2262: out_word = 8'h22;
		16'h2263: out_word = 8'h07;
		16'h2264: out_word = 8'h07;
		16'h2265: out_word = 8'hE6;
		16'h2266: out_word = 8'h50;
		16'h2267: out_word = 8'h47;
		16'h2268: out_word = 8'h3E;
		16'h2269: out_word = 8'h08;
		16'h226A: out_word = 8'hBA;
		16'h226B: out_word = 8'h9F;
		16'h226C: out_word = 8'hAE;
		16'h226D: out_word = 8'hA0;
		16'h226E: out_word = 8'hAE;
		16'h226F: out_word = 8'h77;
		16'h2270: out_word = 8'h23;
		16'h2271: out_word = 8'h78;
		16'h2272: out_word = 8'hC9;
		16'h2273: out_word = 8'h9F;
		16'h2274: out_word = 8'h7A;
		16'h2275: out_word = 8'h0F;
		16'h2276: out_word = 8'h06;
		16'h2277: out_word = 8'h80;
		16'h2278: out_word = 8'h20;
		16'h2279: out_word = 8'h03;
		16'h227A: out_word = 8'h0F;
		16'h227B: out_word = 8'h06;
		16'h227C: out_word = 8'h40;
		16'h227D: out_word = 8'h4F;
		16'h227E: out_word = 8'h7A;
		16'h227F: out_word = 8'hFE;
		16'h2280: out_word = 8'h08;
		16'h2281: out_word = 8'h28;
		16'h2282: out_word = 8'h04;
		16'h2283: out_word = 8'hFE;
		16'h2284: out_word = 8'h02;
		16'h2285: out_word = 8'h30;
		16'h2286: out_word = 8'hBD;
		16'h2287: out_word = 8'h79;
		16'h2288: out_word = 8'h21;
		16'h2289: out_word = 8'h8F;
		16'h228A: out_word = 8'h5C;
		16'h228B: out_word = 8'hCD;
		16'h228C: out_word = 8'h6C;
		16'h228D: out_word = 8'h22;
		16'h228E: out_word = 8'h79;
		16'h228F: out_word = 8'h0F;
		16'h2290: out_word = 8'h0F;
		16'h2291: out_word = 8'h0F;
		16'h2292: out_word = 8'h18;
		16'h2293: out_word = 8'hD8;
		16'h2294: out_word = 8'hCD;
		16'h2295: out_word = 8'h94;
		16'h2296: out_word = 8'h1E;
		16'h2297: out_word = 8'hFE;
		16'h2298: out_word = 8'h08;
		16'h2299: out_word = 8'h30;
		16'h229A: out_word = 8'hA9;
		16'h229B: out_word = 8'hD3;
		16'h229C: out_word = 8'hFE;
		16'h229D: out_word = 8'h07;
		16'h229E: out_word = 8'h07;
		16'h229F: out_word = 8'h07;
		16'h22A0: out_word = 8'hCB;
		16'h22A1: out_word = 8'h6F;
		16'h22A2: out_word = 8'h20;
		16'h22A3: out_word = 8'h02;
		16'h22A4: out_word = 8'hEE;
		16'h22A5: out_word = 8'h07;
		16'h22A6: out_word = 8'h32;
		16'h22A7: out_word = 8'h48;
		16'h22A8: out_word = 8'h5C;
		16'h22A9: out_word = 8'hC9;
		16'h22AA: out_word = 8'h3E;
		16'h22AB: out_word = 8'hAF;
		16'h22AC: out_word = 8'h90;
		16'h22AD: out_word = 8'hDA;
		16'h22AE: out_word = 8'hF9;
		16'h22AF: out_word = 8'h24;
		16'h22B0: out_word = 8'h47;
		16'h22B1: out_word = 8'hA7;
		16'h22B2: out_word = 8'h1F;
		16'h22B3: out_word = 8'h37;
		16'h22B4: out_word = 8'h1F;
		16'h22B5: out_word = 8'hA7;
		16'h22B6: out_word = 8'h1F;
		16'h22B7: out_word = 8'hA8;
		16'h22B8: out_word = 8'hE6;
		16'h22B9: out_word = 8'hF8;
		16'h22BA: out_word = 8'hA8;
		16'h22BB: out_word = 8'h67;
		16'h22BC: out_word = 8'h79;
		16'h22BD: out_word = 8'h07;
		16'h22BE: out_word = 8'h07;
		16'h22BF: out_word = 8'h07;
		16'h22C0: out_word = 8'hA8;
		16'h22C1: out_word = 8'hE6;
		16'h22C2: out_word = 8'hC7;
		16'h22C3: out_word = 8'hA8;
		16'h22C4: out_word = 8'h07;
		16'h22C5: out_word = 8'h07;
		16'h22C6: out_word = 8'h6F;
		16'h22C7: out_word = 8'h79;
		16'h22C8: out_word = 8'hE6;
		16'h22C9: out_word = 8'h07;
		16'h22CA: out_word = 8'hC9;
		16'h22CB: out_word = 8'hCD;
		16'h22CC: out_word = 8'h07;
		16'h22CD: out_word = 8'h23;
		16'h22CE: out_word = 8'hCD;
		16'h22CF: out_word = 8'hAA;
		16'h22D0: out_word = 8'h22;
		16'h22D1: out_word = 8'h47;
		16'h22D2: out_word = 8'h04;
		16'h22D3: out_word = 8'h7E;
		16'h22D4: out_word = 8'h07;
		16'h22D5: out_word = 8'h10;
		16'h22D6: out_word = 8'hFD;
		16'h22D7: out_word = 8'hE6;
		16'h22D8: out_word = 8'h01;
		16'h22D9: out_word = 8'hC3;
		16'h22DA: out_word = 8'h28;
		16'h22DB: out_word = 8'h2D;
		16'h22DC: out_word = 8'hCD;
		16'h22DD: out_word = 8'h07;
		16'h22DE: out_word = 8'h23;
		16'h22DF: out_word = 8'hCD;
		16'h22E0: out_word = 8'hE5;
		16'h22E1: out_word = 8'h22;
		16'h22E2: out_word = 8'hC3;
		16'h22E3: out_word = 8'h4D;
		16'h22E4: out_word = 8'h0D;
		16'h22E5: out_word = 8'hED;
		16'h22E6: out_word = 8'h43;
		16'h22E7: out_word = 8'h7D;
		16'h22E8: out_word = 8'h5C;
		16'h22E9: out_word = 8'hCD;
		16'h22EA: out_word = 8'hAA;
		16'h22EB: out_word = 8'h22;
		16'h22EC: out_word = 8'h47;
		16'h22ED: out_word = 8'h04;
		16'h22EE: out_word = 8'h3E;
		16'h22EF: out_word = 8'hFE;
		16'h22F0: out_word = 8'h0F;
		16'h22F1: out_word = 8'h10;
		16'h22F2: out_word = 8'hFD;
		16'h22F3: out_word = 8'h47;
		16'h22F4: out_word = 8'h7E;
		16'h22F5: out_word = 8'hFD;
		16'h22F6: out_word = 8'h4E;
		16'h22F7: out_word = 8'h57;
		16'h22F8: out_word = 8'hCB;
		16'h22F9: out_word = 8'h41;
		16'h22FA: out_word = 8'h20;
		16'h22FB: out_word = 8'h01;
		16'h22FC: out_word = 8'hA0;
		16'h22FD: out_word = 8'hCB;
		16'h22FE: out_word = 8'h51;
		16'h22FF: out_word = 8'h20;
		16'h2300: out_word = 8'h02;
		16'h2301: out_word = 8'hA8;
		16'h2302: out_word = 8'h2F;
		16'h2303: out_word = 8'h77;
		16'h2304: out_word = 8'hC3;
		16'h2305: out_word = 8'hDB;
		16'h2306: out_word = 8'h0B;
		16'h2307: out_word = 8'hCD;
		16'h2308: out_word = 8'h14;
		16'h2309: out_word = 8'h23;
		16'h230A: out_word = 8'h47;
		16'h230B: out_word = 8'hC5;
		16'h230C: out_word = 8'hCD;
		16'h230D: out_word = 8'h14;
		16'h230E: out_word = 8'h23;
		16'h230F: out_word = 8'h59;
		16'h2310: out_word = 8'hC1;
		16'h2311: out_word = 8'h51;
		16'h2312: out_word = 8'h4F;
		16'h2313: out_word = 8'hC9;
		16'h2314: out_word = 8'hCD;
		16'h2315: out_word = 8'hD5;
		16'h2316: out_word = 8'h2D;
		16'h2317: out_word = 8'hDA;
		16'h2318: out_word = 8'hF9;
		16'h2319: out_word = 8'h24;
		16'h231A: out_word = 8'h0E;
		16'h231B: out_word = 8'h01;
		16'h231C: out_word = 8'hC8;
		16'h231D: out_word = 8'h0E;
		16'h231E: out_word = 8'hFF;
		16'h231F: out_word = 8'hC9;
		16'h2320: out_word = 8'hDF;
		16'h2321: out_word = 8'hFE;
		16'h2322: out_word = 8'h2C;
		16'h2323: out_word = 8'hC2;
		16'h2324: out_word = 8'h8A;
		16'h2325: out_word = 8'h1C;
		16'h2326: out_word = 8'hE7;
		16'h2327: out_word = 8'hCD;
		16'h2328: out_word = 8'h82;
		16'h2329: out_word = 8'h1C;
		16'h232A: out_word = 8'hCD;
		16'h232B: out_word = 8'hEE;
		16'h232C: out_word = 8'h1B;
		16'h232D: out_word = 8'hEF;
		16'h232E: out_word = 8'h2A;
		16'h232F: out_word = 8'h3D;
		16'h2330: out_word = 8'h38;
		16'h2331: out_word = 8'h7E;
		16'h2332: out_word = 8'hFE;
		16'h2333: out_word = 8'h81;
		16'h2334: out_word = 8'h30;
		16'h2335: out_word = 8'h05;
		16'h2336: out_word = 8'hEF;
		16'h2337: out_word = 8'h02;
		16'h2338: out_word = 8'h38;
		16'h2339: out_word = 8'h18;
		16'h233A: out_word = 8'hA1;
		16'h233B: out_word = 8'hEF;
		16'h233C: out_word = 8'hA3;
		16'h233D: out_word = 8'h38;
		16'h233E: out_word = 8'h36;
		16'h233F: out_word = 8'h83;
		16'h2340: out_word = 8'hEF;
		16'h2341: out_word = 8'hC5;
		16'h2342: out_word = 8'h02;
		16'h2343: out_word = 8'h38;
		16'h2344: out_word = 8'hCD;
		16'h2345: out_word = 8'h7D;
		16'h2346: out_word = 8'h24;
		16'h2347: out_word = 8'hC5;
		16'h2348: out_word = 8'hEF;
		16'h2349: out_word = 8'h31;
		16'h234A: out_word = 8'hE1;
		16'h234B: out_word = 8'h04;
		16'h234C: out_word = 8'h38;
		16'h234D: out_word = 8'h7E;
		16'h234E: out_word = 8'hFE;
		16'h234F: out_word = 8'h80;
		16'h2350: out_word = 8'h30;
		16'h2351: out_word = 8'h08;
		16'h2352: out_word = 8'hEF;
		16'h2353: out_word = 8'h02;
		16'h2354: out_word = 8'h02;
		16'h2355: out_word = 8'h38;
		16'h2356: out_word = 8'hC1;
		16'h2357: out_word = 8'hC3;
		16'h2358: out_word = 8'hDC;
		16'h2359: out_word = 8'h22;
		16'h235A: out_word = 8'hEF;
		16'h235B: out_word = 8'hC2;
		16'h235C: out_word = 8'h01;
		16'h235D: out_word = 8'hC0;
		16'h235E: out_word = 8'h02;
		16'h235F: out_word = 8'h03;
		16'h2360: out_word = 8'h01;
		16'h2361: out_word = 8'hE0;
		16'h2362: out_word = 8'h0F;
		16'h2363: out_word = 8'hC0;
		16'h2364: out_word = 8'h01;
		16'h2365: out_word = 8'h31;
		16'h2366: out_word = 8'hE0;
		16'h2367: out_word = 8'h01;
		16'h2368: out_word = 8'h31;
		16'h2369: out_word = 8'hE0;
		16'h236A: out_word = 8'hA0;
		16'h236B: out_word = 8'hC1;
		16'h236C: out_word = 8'h02;
		16'h236D: out_word = 8'h38;
		16'h236E: out_word = 8'hFD;
		16'h236F: out_word = 8'h34;
		16'h2370: out_word = 8'h62;
		16'h2371: out_word = 8'hCD;
		16'h2372: out_word = 8'h94;
		16'h2373: out_word = 8'h1E;
		16'h2374: out_word = 8'h6F;
		16'h2375: out_word = 8'hE5;
		16'h2376: out_word = 8'hCD;
		16'h2377: out_word = 8'h94;
		16'h2378: out_word = 8'h1E;
		16'h2379: out_word = 8'hE1;
		16'h237A: out_word = 8'h67;
		16'h237B: out_word = 8'h22;
		16'h237C: out_word = 8'h7D;
		16'h237D: out_word = 8'h5C;
		16'h237E: out_word = 8'hC1;
		16'h237F: out_word = 8'hC3;
		16'h2380: out_word = 8'h20;
		16'h2381: out_word = 8'h24;
		16'h2382: out_word = 8'hDF;
		16'h2383: out_word = 8'hFE;
		16'h2384: out_word = 8'h2C;
		16'h2385: out_word = 8'h28;
		16'h2386: out_word = 8'h06;
		16'h2387: out_word = 8'hCD;
		16'h2388: out_word = 8'hEE;
		16'h2389: out_word = 8'h1B;
		16'h238A: out_word = 8'hC3;
		16'h238B: out_word = 8'h77;
		16'h238C: out_word = 8'h24;
		16'h238D: out_word = 8'hE7;
		16'h238E: out_word = 8'hCD;
		16'h238F: out_word = 8'h82;
		16'h2390: out_word = 8'h1C;
		16'h2391: out_word = 8'hCD;
		16'h2392: out_word = 8'hEE;
		16'h2393: out_word = 8'h1B;
		16'h2394: out_word = 8'hEF;
		16'h2395: out_word = 8'hC5;
		16'h2396: out_word = 8'hA2;
		16'h2397: out_word = 8'h04;
		16'h2398: out_word = 8'h1F;
		16'h2399: out_word = 8'h31;
		16'h239A: out_word = 8'h30;
		16'h239B: out_word = 8'h30;
		16'h239C: out_word = 8'h00;
		16'h239D: out_word = 8'h06;
		16'h239E: out_word = 8'h02;
		16'h239F: out_word = 8'h38;
		16'h23A0: out_word = 8'hC3;
		16'h23A1: out_word = 8'h77;
		16'h23A2: out_word = 8'h24;
		16'h23A3: out_word = 8'hC0;
		16'h23A4: out_word = 8'h02;
		16'h23A5: out_word = 8'hC1;
		16'h23A6: out_word = 8'h02;
		16'h23A7: out_word = 8'h31;
		16'h23A8: out_word = 8'h2A;
		16'h23A9: out_word = 8'hE1;
		16'h23AA: out_word = 8'h01;
		16'h23AB: out_word = 8'hE1;
		16'h23AC: out_word = 8'h2A;
		16'h23AD: out_word = 8'h0F;
		16'h23AE: out_word = 8'hE0;
		16'h23AF: out_word = 8'h05;
		16'h23B0: out_word = 8'h2A;
		16'h23B1: out_word = 8'hE0;
		16'h23B2: out_word = 8'h01;
		16'h23B3: out_word = 8'h3D;
		16'h23B4: out_word = 8'h38;
		16'h23B5: out_word = 8'h7E;
		16'h23B6: out_word = 8'hFE;
		16'h23B7: out_word = 8'h81;
		16'h23B8: out_word = 8'h30;
		16'h23B9: out_word = 8'h07;
		16'h23BA: out_word = 8'hEF;
		16'h23BB: out_word = 8'h02;
		16'h23BC: out_word = 8'h02;
		16'h23BD: out_word = 8'h38;
		16'h23BE: out_word = 8'hC3;
		16'h23BF: out_word = 8'h77;
		16'h23C0: out_word = 8'h24;
		16'h23C1: out_word = 8'hCD;
		16'h23C2: out_word = 8'h7D;
		16'h23C3: out_word = 8'h24;
		16'h23C4: out_word = 8'hC5;
		16'h23C5: out_word = 8'hEF;
		16'h23C6: out_word = 8'h02;
		16'h23C7: out_word = 8'hE1;
		16'h23C8: out_word = 8'h01;
		16'h23C9: out_word = 8'h05;
		16'h23CA: out_word = 8'hC1;
		16'h23CB: out_word = 8'h02;
		16'h23CC: out_word = 8'h01;
		16'h23CD: out_word = 8'h31;
		16'h23CE: out_word = 8'hE1;
		16'h23CF: out_word = 8'h04;
		16'h23D0: out_word = 8'hC2;
		16'h23D1: out_word = 8'h02;
		16'h23D2: out_word = 8'h01;
		16'h23D3: out_word = 8'h31;
		16'h23D4: out_word = 8'hE1;
		16'h23D5: out_word = 8'h04;
		16'h23D6: out_word = 8'hE2;
		16'h23D7: out_word = 8'hE5;
		16'h23D8: out_word = 8'hE0;
		16'h23D9: out_word = 8'h03;
		16'h23DA: out_word = 8'hA2;
		16'h23DB: out_word = 8'h04;
		16'h23DC: out_word = 8'h31;
		16'h23DD: out_word = 8'h1F;
		16'h23DE: out_word = 8'hC5;
		16'h23DF: out_word = 8'h02;
		16'h23E0: out_word = 8'h20;
		16'h23E1: out_word = 8'hC0;
		16'h23E2: out_word = 8'h02;
		16'h23E3: out_word = 8'hC2;
		16'h23E4: out_word = 8'h02;
		16'h23E5: out_word = 8'hC1;
		16'h23E6: out_word = 8'hE5;
		16'h23E7: out_word = 8'h04;
		16'h23E8: out_word = 8'hE0;
		16'h23E9: out_word = 8'hE2;
		16'h23EA: out_word = 8'h04;
		16'h23EB: out_word = 8'h0F;
		16'h23EC: out_word = 8'hE1;
		16'h23ED: out_word = 8'h01;
		16'h23EE: out_word = 8'hC1;
		16'h23EF: out_word = 8'h02;
		16'h23F0: out_word = 8'hE0;
		16'h23F1: out_word = 8'h04;
		16'h23F2: out_word = 8'hE2;
		16'h23F3: out_word = 8'hE5;
		16'h23F4: out_word = 8'h04;
		16'h23F5: out_word = 8'h03;
		16'h23F6: out_word = 8'hC2;
		16'h23F7: out_word = 8'h2A;
		16'h23F8: out_word = 8'hE1;
		16'h23F9: out_word = 8'h2A;
		16'h23FA: out_word = 8'h0F;
		16'h23FB: out_word = 8'h02;
		16'h23FC: out_word = 8'h38;
		16'h23FD: out_word = 8'h1A;
		16'h23FE: out_word = 8'hFE;
		16'h23FF: out_word = 8'h81;
		16'h2400: out_word = 8'hC1;
		16'h2401: out_word = 8'hDA;
		16'h2402: out_word = 8'h77;
		16'h2403: out_word = 8'h24;
		16'h2404: out_word = 8'hC5;
		16'h2405: out_word = 8'hEF;
		16'h2406: out_word = 8'h01;
		16'h2407: out_word = 8'h38;
		16'h2408: out_word = 8'h3A;
		16'h2409: out_word = 8'h7D;
		16'h240A: out_word = 8'h5C;
		16'h240B: out_word = 8'hCD;
		16'h240C: out_word = 8'h28;
		16'h240D: out_word = 8'h2D;
		16'h240E: out_word = 8'hEF;
		16'h240F: out_word = 8'hC0;
		16'h2410: out_word = 8'h0F;
		16'h2411: out_word = 8'h01;
		16'h2412: out_word = 8'h38;
		16'h2413: out_word = 8'h3A;
		16'h2414: out_word = 8'h7E;
		16'h2415: out_word = 8'h5C;
		16'h2416: out_word = 8'hCD;
		16'h2417: out_word = 8'h28;
		16'h2418: out_word = 8'h2D;
		16'h2419: out_word = 8'hEF;
		16'h241A: out_word = 8'hC5;
		16'h241B: out_word = 8'h0F;
		16'h241C: out_word = 8'hE0;
		16'h241D: out_word = 8'hE5;
		16'h241E: out_word = 8'h38;
		16'h241F: out_word = 8'hC1;
		16'h2420: out_word = 8'h05;
		16'h2421: out_word = 8'h28;
		16'h2422: out_word = 8'h3C;
		16'h2423: out_word = 8'h18;
		16'h2424: out_word = 8'h14;
		16'h2425: out_word = 8'hEF;
		16'h2426: out_word = 8'hE1;
		16'h2427: out_word = 8'h31;
		16'h2428: out_word = 8'hE3;
		16'h2429: out_word = 8'h04;
		16'h242A: out_word = 8'hE2;
		16'h242B: out_word = 8'hE4;
		16'h242C: out_word = 8'h04;
		16'h242D: out_word = 8'h03;
		16'h242E: out_word = 8'hC1;
		16'h242F: out_word = 8'h02;
		16'h2430: out_word = 8'hE4;
		16'h2431: out_word = 8'h04;
		16'h2432: out_word = 8'hE2;
		16'h2433: out_word = 8'hE3;
		16'h2434: out_word = 8'h04;
		16'h2435: out_word = 8'h0F;
		16'h2436: out_word = 8'hC2;
		16'h2437: out_word = 8'h02;
		16'h2438: out_word = 8'h38;
		16'h2439: out_word = 8'hC5;
		16'h243A: out_word = 8'hEF;
		16'h243B: out_word = 8'hC0;
		16'h243C: out_word = 8'h02;
		16'h243D: out_word = 8'hE1;
		16'h243E: out_word = 8'h0F;
		16'h243F: out_word = 8'h31;
		16'h2440: out_word = 8'h38;
		16'h2441: out_word = 8'h3A;
		16'h2442: out_word = 8'h7D;
		16'h2443: out_word = 8'h5C;
		16'h2444: out_word = 8'hCD;
		16'h2445: out_word = 8'h28;
		16'h2446: out_word = 8'h2D;
		16'h2447: out_word = 8'hEF;
		16'h2448: out_word = 8'h03;
		16'h2449: out_word = 8'hE0;
		16'h244A: out_word = 8'hE2;
		16'h244B: out_word = 8'h0F;
		16'h244C: out_word = 8'hC0;
		16'h244D: out_word = 8'h01;
		16'h244E: out_word = 8'hE0;
		16'h244F: out_word = 8'h38;
		16'h2450: out_word = 8'h3A;
		16'h2451: out_word = 8'h7E;
		16'h2452: out_word = 8'h5C;
		16'h2453: out_word = 8'hCD;
		16'h2454: out_word = 8'h28;
		16'h2455: out_word = 8'h2D;
		16'h2456: out_word = 8'hEF;
		16'h2457: out_word = 8'h03;
		16'h2458: out_word = 8'h38;
		16'h2459: out_word = 8'hCD;
		16'h245A: out_word = 8'hB7;
		16'h245B: out_word = 8'h24;
		16'h245C: out_word = 8'hC1;
		16'h245D: out_word = 8'h10;
		16'h245E: out_word = 8'hC6;
		16'h245F: out_word = 8'hEF;
		16'h2460: out_word = 8'h02;
		16'h2461: out_word = 8'h02;
		16'h2462: out_word = 8'h01;
		16'h2463: out_word = 8'h38;
		16'h2464: out_word = 8'h3A;
		16'h2465: out_word = 8'h7D;
		16'h2466: out_word = 8'h5C;
		16'h2467: out_word = 8'hCD;
		16'h2468: out_word = 8'h28;
		16'h2469: out_word = 8'h2D;
		16'h246A: out_word = 8'hEF;
		16'h246B: out_word = 8'h03;
		16'h246C: out_word = 8'h01;
		16'h246D: out_word = 8'h38;
		16'h246E: out_word = 8'h3A;
		16'h246F: out_word = 8'h7E;
		16'h2470: out_word = 8'h5C;
		16'h2471: out_word = 8'hCD;
		16'h2472: out_word = 8'h28;
		16'h2473: out_word = 8'h2D;
		16'h2474: out_word = 8'hEF;
		16'h2475: out_word = 8'h03;
		16'h2476: out_word = 8'h38;
		16'h2477: out_word = 8'hCD;
		16'h2478: out_word = 8'hB7;
		16'h2479: out_word = 8'h24;
		16'h247A: out_word = 8'hC3;
		16'h247B: out_word = 8'h4D;
		16'h247C: out_word = 8'h0D;
		16'h247D: out_word = 8'hEF;
		16'h247E: out_word = 8'h31;
		16'h247F: out_word = 8'h28;
		16'h2480: out_word = 8'h34;
		16'h2481: out_word = 8'h32;
		16'h2482: out_word = 8'h00;
		16'h2483: out_word = 8'h01;
		16'h2484: out_word = 8'h05;
		16'h2485: out_word = 8'hE5;
		16'h2486: out_word = 8'h01;
		16'h2487: out_word = 8'h05;
		16'h2488: out_word = 8'h2A;
		16'h2489: out_word = 8'h38;
		16'h248A: out_word = 8'hCD;
		16'h248B: out_word = 8'hD5;
		16'h248C: out_word = 8'h2D;
		16'h248D: out_word = 8'h38;
		16'h248E: out_word = 8'h06;
		16'h248F: out_word = 8'hE6;
		16'h2490: out_word = 8'hFC;
		16'h2491: out_word = 8'hC6;
		16'h2492: out_word = 8'h04;
		16'h2493: out_word = 8'h30;
		16'h2494: out_word = 8'h02;
		16'h2495: out_word = 8'h3E;
		16'h2496: out_word = 8'hFC;
		16'h2497: out_word = 8'hF5;
		16'h2498: out_word = 8'hCD;
		16'h2499: out_word = 8'h28;
		16'h249A: out_word = 8'h2D;
		16'h249B: out_word = 8'hEF;
		16'h249C: out_word = 8'hE5;
		16'h249D: out_word = 8'h01;
		16'h249E: out_word = 8'h05;
		16'h249F: out_word = 8'h31;
		16'h24A0: out_word = 8'h1F;
		16'h24A1: out_word = 8'hC4;
		16'h24A2: out_word = 8'h02;
		16'h24A3: out_word = 8'h31;
		16'h24A4: out_word = 8'hA2;
		16'h24A5: out_word = 8'h04;
		16'h24A6: out_word = 8'h1F;
		16'h24A7: out_word = 8'hC1;
		16'h24A8: out_word = 8'h01;
		16'h24A9: out_word = 8'hC0;
		16'h24AA: out_word = 8'h02;
		16'h24AB: out_word = 8'h31;
		16'h24AC: out_word = 8'h04;
		16'h24AD: out_word = 8'h31;
		16'h24AE: out_word = 8'h0F;
		16'h24AF: out_word = 8'hA1;
		16'h24B0: out_word = 8'h03;
		16'h24B1: out_word = 8'h1B;
		16'h24B2: out_word = 8'hC3;
		16'h24B3: out_word = 8'h02;
		16'h24B4: out_word = 8'h38;
		16'h24B5: out_word = 8'hC1;
		16'h24B6: out_word = 8'hC9;
		16'h24B7: out_word = 8'hCD;
		16'h24B8: out_word = 8'h07;
		16'h24B9: out_word = 8'h23;
		16'h24BA: out_word = 8'h79;
		16'h24BB: out_word = 8'hB8;
		16'h24BC: out_word = 8'h30;
		16'h24BD: out_word = 8'h06;
		16'h24BE: out_word = 8'h69;
		16'h24BF: out_word = 8'hD5;
		16'h24C0: out_word = 8'hAF;
		16'h24C1: out_word = 8'h5F;
		16'h24C2: out_word = 8'h18;
		16'h24C3: out_word = 8'h07;
		16'h24C4: out_word = 8'hB1;
		16'h24C5: out_word = 8'hC8;
		16'h24C6: out_word = 8'h68;
		16'h24C7: out_word = 8'h41;
		16'h24C8: out_word = 8'hD5;
		16'h24C9: out_word = 8'h16;
		16'h24CA: out_word = 8'h00;
		16'h24CB: out_word = 8'h60;
		16'h24CC: out_word = 8'h78;
		16'h24CD: out_word = 8'h1F;
		16'h24CE: out_word = 8'h85;
		16'h24CF: out_word = 8'h38;
		16'h24D0: out_word = 8'h03;
		16'h24D1: out_word = 8'hBC;
		16'h24D2: out_word = 8'h38;
		16'h24D3: out_word = 8'h07;
		16'h24D4: out_word = 8'h94;
		16'h24D5: out_word = 8'h4F;
		16'h24D6: out_word = 8'hD9;
		16'h24D7: out_word = 8'hC1;
		16'h24D8: out_word = 8'hC5;
		16'h24D9: out_word = 8'h18;
		16'h24DA: out_word = 8'h04;
		16'h24DB: out_word = 8'h4F;
		16'h24DC: out_word = 8'hD5;
		16'h24DD: out_word = 8'hD9;
		16'h24DE: out_word = 8'hC1;
		16'h24DF: out_word = 8'h2A;
		16'h24E0: out_word = 8'h7D;
		16'h24E1: out_word = 8'h5C;
		16'h24E2: out_word = 8'h78;
		16'h24E3: out_word = 8'h84;
		16'h24E4: out_word = 8'h47;
		16'h24E5: out_word = 8'h79;
		16'h24E6: out_word = 8'h3C;
		16'h24E7: out_word = 8'h85;
		16'h24E8: out_word = 8'h38;
		16'h24E9: out_word = 8'h0D;
		16'h24EA: out_word = 8'h28;
		16'h24EB: out_word = 8'h0D;
		16'h24EC: out_word = 8'h3D;
		16'h24ED: out_word = 8'h4F;
		16'h24EE: out_word = 8'hCD;
		16'h24EF: out_word = 8'hE5;
		16'h24F0: out_word = 8'h22;
		16'h24F1: out_word = 8'hD9;
		16'h24F2: out_word = 8'h79;
		16'h24F3: out_word = 8'h10;
		16'h24F4: out_word = 8'hD9;
		16'h24F5: out_word = 8'hD1;
		16'h24F6: out_word = 8'hC9;
		16'h24F7: out_word = 8'h28;
		16'h24F8: out_word = 8'hF3;
		16'h24F9: out_word = 8'hCF;
		16'h24FA: out_word = 8'h0A;
		16'h24FB: out_word = 8'hDF;
		16'h24FC: out_word = 8'h06;
		16'h24FD: out_word = 8'h00;
		16'h24FE: out_word = 8'hC5;
		16'h24FF: out_word = 8'h4F;
		16'h2500: out_word = 8'h21;
		16'h2501: out_word = 8'h96;
		16'h2502: out_word = 8'h25;
		16'h2503: out_word = 8'hCD;
		16'h2504: out_word = 8'hDC;
		16'h2505: out_word = 8'h16;
		16'h2506: out_word = 8'h79;
		16'h2507: out_word = 8'hD2;
		16'h2508: out_word = 8'h84;
		16'h2509: out_word = 8'h26;
		16'h250A: out_word = 8'h06;
		16'h250B: out_word = 8'h00;
		16'h250C: out_word = 8'h4E;
		16'h250D: out_word = 8'h09;
		16'h250E: out_word = 8'hE9;
		16'h250F: out_word = 8'hCD;
		16'h2510: out_word = 8'h74;
		16'h2511: out_word = 8'h00;
		16'h2512: out_word = 8'h03;
		16'h2513: out_word = 8'hFE;
		16'h2514: out_word = 8'h0D;
		16'h2515: out_word = 8'hCA;
		16'h2516: out_word = 8'h8A;
		16'h2517: out_word = 8'h1C;
		16'h2518: out_word = 8'hFE;
		16'h2519: out_word = 8'h22;
		16'h251A: out_word = 8'h20;
		16'h251B: out_word = 8'hF3;
		16'h251C: out_word = 8'hCD;
		16'h251D: out_word = 8'h74;
		16'h251E: out_word = 8'h00;
		16'h251F: out_word = 8'hFE;
		16'h2520: out_word = 8'h22;
		16'h2521: out_word = 8'hC9;
		16'h2522: out_word = 8'hE7;
		16'h2523: out_word = 8'hFE;
		16'h2524: out_word = 8'h28;
		16'h2525: out_word = 8'h20;
		16'h2526: out_word = 8'h06;
		16'h2527: out_word = 8'hCD;
		16'h2528: out_word = 8'h79;
		16'h2529: out_word = 8'h1C;
		16'h252A: out_word = 8'hDF;
		16'h252B: out_word = 8'hFE;
		16'h252C: out_word = 8'h29;
		16'h252D: out_word = 8'hC2;
		16'h252E: out_word = 8'h8A;
		16'h252F: out_word = 8'h1C;
		16'h2530: out_word = 8'hFD;
		16'h2531: out_word = 8'hCB;
		16'h2532: out_word = 8'h01;
		16'h2533: out_word = 8'h7E;
		16'h2534: out_word = 8'hC9;
		16'h2535: out_word = 8'hCD;
		16'h2536: out_word = 8'h07;
		16'h2537: out_word = 8'h23;
		16'h2538: out_word = 8'h2A;
		16'h2539: out_word = 8'h36;
		16'h253A: out_word = 8'h5C;
		16'h253B: out_word = 8'h11;
		16'h253C: out_word = 8'h00;
		16'h253D: out_word = 8'h01;
		16'h253E: out_word = 8'h19;
		16'h253F: out_word = 8'h79;
		16'h2540: out_word = 8'h0F;
		16'h2541: out_word = 8'h0F;
		16'h2542: out_word = 8'h0F;
		16'h2543: out_word = 8'hE6;
		16'h2544: out_word = 8'hE0;
		16'h2545: out_word = 8'hA8;
		16'h2546: out_word = 8'h5F;
		16'h2547: out_word = 8'h79;
		16'h2548: out_word = 8'hE6;
		16'h2549: out_word = 8'h18;
		16'h254A: out_word = 8'hEE;
		16'h254B: out_word = 8'h40;
		16'h254C: out_word = 8'h57;
		16'h254D: out_word = 8'h06;
		16'h254E: out_word = 8'h60;
		16'h254F: out_word = 8'hC5;
		16'h2550: out_word = 8'hD5;
		16'h2551: out_word = 8'hE5;
		16'h2552: out_word = 8'h1A;
		16'h2553: out_word = 8'hAE;
		16'h2554: out_word = 8'h28;
		16'h2555: out_word = 8'h04;
		16'h2556: out_word = 8'h3C;
		16'h2557: out_word = 8'h20;
		16'h2558: out_word = 8'h1A;
		16'h2559: out_word = 8'h3D;
		16'h255A: out_word = 8'h4F;
		16'h255B: out_word = 8'h06;
		16'h255C: out_word = 8'h07;
		16'h255D: out_word = 8'h14;
		16'h255E: out_word = 8'h23;
		16'h255F: out_word = 8'h1A;
		16'h2560: out_word = 8'hAE;
		16'h2561: out_word = 8'hA9;
		16'h2562: out_word = 8'h20;
		16'h2563: out_word = 8'h0F;
		16'h2564: out_word = 8'h10;
		16'h2565: out_word = 8'hF7;
		16'h2566: out_word = 8'hC1;
		16'h2567: out_word = 8'hC1;
		16'h2568: out_word = 8'hC1;
		16'h2569: out_word = 8'h3E;
		16'h256A: out_word = 8'h80;
		16'h256B: out_word = 8'h90;
		16'h256C: out_word = 8'h01;
		16'h256D: out_word = 8'h01;
		16'h256E: out_word = 8'h00;
		16'h256F: out_word = 8'hF7;
		16'h2570: out_word = 8'h12;
		16'h2571: out_word = 8'h18;
		16'h2572: out_word = 8'h0A;
		16'h2573: out_word = 8'hE1;
		16'h2574: out_word = 8'h11;
		16'h2575: out_word = 8'h08;
		16'h2576: out_word = 8'h00;
		16'h2577: out_word = 8'h19;
		16'h2578: out_word = 8'hD1;
		16'h2579: out_word = 8'hC1;
		16'h257A: out_word = 8'h10;
		16'h257B: out_word = 8'hD3;
		16'h257C: out_word = 8'h48;
		16'h257D: out_word = 8'hC3;
		16'h257E: out_word = 8'hB2;
		16'h257F: out_word = 8'h2A;
		16'h2580: out_word = 8'hCD;
		16'h2581: out_word = 8'h07;
		16'h2582: out_word = 8'h23;
		16'h2583: out_word = 8'h79;
		16'h2584: out_word = 8'h0F;
		16'h2585: out_word = 8'h0F;
		16'h2586: out_word = 8'h0F;
		16'h2587: out_word = 8'h4F;
		16'h2588: out_word = 8'hE6;
		16'h2589: out_word = 8'hE0;
		16'h258A: out_word = 8'hA8;
		16'h258B: out_word = 8'h6F;
		16'h258C: out_word = 8'h79;
		16'h258D: out_word = 8'hE6;
		16'h258E: out_word = 8'h03;
		16'h258F: out_word = 8'hEE;
		16'h2590: out_word = 8'h58;
		16'h2591: out_word = 8'h67;
		16'h2592: out_word = 8'h7E;
		16'h2593: out_word = 8'hC3;
		16'h2594: out_word = 8'h28;
		16'h2595: out_word = 8'h2D;
		16'h2596: out_word = 8'h22;
		16'h2597: out_word = 8'h1C;
		16'h2598: out_word = 8'h28;
		16'h2599: out_word = 8'h4F;
		16'h259A: out_word = 8'h2E;
		16'h259B: out_word = 8'hF2;
		16'h259C: out_word = 8'h2B;
		16'h259D: out_word = 8'h12;
		16'h259E: out_word = 8'hA8;
		16'h259F: out_word = 8'h56;
		16'h25A0: out_word = 8'hA5;
		16'h25A1: out_word = 8'h57;
		16'h25A2: out_word = 8'hA7;
		16'h25A3: out_word = 8'h84;
		16'h25A4: out_word = 8'hA6;
		16'h25A5: out_word = 8'h8F;
		16'h25A6: out_word = 8'hC4;
		16'h25A7: out_word = 8'hE6;
		16'h25A8: out_word = 8'hAA;
		16'h25A9: out_word = 8'hBF;
		16'h25AA: out_word = 8'hAB;
		16'h25AB: out_word = 8'hC7;
		16'h25AC: out_word = 8'hA9;
		16'h25AD: out_word = 8'hCE;
		16'h25AE: out_word = 8'h00;
		16'h25AF: out_word = 8'hE7;
		16'h25B0: out_word = 8'hC3;
		16'h25B1: out_word = 8'hFF;
		16'h25B2: out_word = 8'h24;
		16'h25B3: out_word = 8'hDF;
		16'h25B4: out_word = 8'h23;
		16'h25B5: out_word = 8'hE5;
		16'h25B6: out_word = 8'h01;
		16'h25B7: out_word = 8'h00;
		16'h25B8: out_word = 8'h00;
		16'h25B9: out_word = 8'hCD;
		16'h25BA: out_word = 8'h0F;
		16'h25BB: out_word = 8'h25;
		16'h25BC: out_word = 8'h20;
		16'h25BD: out_word = 8'h1B;
		16'h25BE: out_word = 8'hCD;
		16'h25BF: out_word = 8'h0F;
		16'h25C0: out_word = 8'h25;
		16'h25C1: out_word = 8'h28;
		16'h25C2: out_word = 8'hFB;
		16'h25C3: out_word = 8'hCD;
		16'h25C4: out_word = 8'h30;
		16'h25C5: out_word = 8'h25;
		16'h25C6: out_word = 8'h28;
		16'h25C7: out_word = 8'h11;
		16'h25C8: out_word = 8'hF7;
		16'h25C9: out_word = 8'hE1;
		16'h25CA: out_word = 8'hD5;
		16'h25CB: out_word = 8'h7E;
		16'h25CC: out_word = 8'h23;
		16'h25CD: out_word = 8'h12;
		16'h25CE: out_word = 8'h13;
		16'h25CF: out_word = 8'hFE;
		16'h25D0: out_word = 8'h22;
		16'h25D1: out_word = 8'h20;
		16'h25D2: out_word = 8'hF8;
		16'h25D3: out_word = 8'h7E;
		16'h25D4: out_word = 8'h23;
		16'h25D5: out_word = 8'hFE;
		16'h25D6: out_word = 8'h22;
		16'h25D7: out_word = 8'h28;
		16'h25D8: out_word = 8'hF2;
		16'h25D9: out_word = 8'h0B;
		16'h25DA: out_word = 8'hD1;
		16'h25DB: out_word = 8'h21;
		16'h25DC: out_word = 8'h3B;
		16'h25DD: out_word = 8'h5C;
		16'h25DE: out_word = 8'hCB;
		16'h25DF: out_word = 8'hB6;
		16'h25E0: out_word = 8'hCB;
		16'h25E1: out_word = 8'h7E;
		16'h25E2: out_word = 8'hC4;
		16'h25E3: out_word = 8'hB2;
		16'h25E4: out_word = 8'h2A;
		16'h25E5: out_word = 8'hC3;
		16'h25E6: out_word = 8'h12;
		16'h25E7: out_word = 8'h27;
		16'h25E8: out_word = 8'hE7;
		16'h25E9: out_word = 8'hCD;
		16'h25EA: out_word = 8'hFB;
		16'h25EB: out_word = 8'h24;
		16'h25EC: out_word = 8'hFE;
		16'h25ED: out_word = 8'h29;
		16'h25EE: out_word = 8'hC2;
		16'h25EF: out_word = 8'h8A;
		16'h25F0: out_word = 8'h1C;
		16'h25F1: out_word = 8'hE7;
		16'h25F2: out_word = 8'hC3;
		16'h25F3: out_word = 8'h12;
		16'h25F4: out_word = 8'h27;
		16'h25F5: out_word = 8'hC3;
		16'h25F6: out_word = 8'hBD;
		16'h25F7: out_word = 8'h27;
		16'h25F8: out_word = 8'hCD;
		16'h25F9: out_word = 8'h30;
		16'h25FA: out_word = 8'h25;
		16'h25FB: out_word = 8'h28;
		16'h25FC: out_word = 8'h28;
		16'h25FD: out_word = 8'hED;
		16'h25FE: out_word = 8'h4B;
		16'h25FF: out_word = 8'h76;
		16'h2600: out_word = 8'h5C;
		16'h2601: out_word = 8'hCD;
		16'h2602: out_word = 8'h2B;
		16'h2603: out_word = 8'h2D;
		16'h2604: out_word = 8'hEF;
		16'h2605: out_word = 8'hA1;
		16'h2606: out_word = 8'h0F;
		16'h2607: out_word = 8'h34;
		16'h2608: out_word = 8'h37;
		16'h2609: out_word = 8'h16;
		16'h260A: out_word = 8'h04;
		16'h260B: out_word = 8'h34;
		16'h260C: out_word = 8'h80;
		16'h260D: out_word = 8'h41;
		16'h260E: out_word = 8'h00;
		16'h260F: out_word = 8'h00;
		16'h2610: out_word = 8'h80;
		16'h2611: out_word = 8'h32;
		16'h2612: out_word = 8'h02;
		16'h2613: out_word = 8'hA1;
		16'h2614: out_word = 8'h03;
		16'h2615: out_word = 8'h31;
		16'h2616: out_word = 8'h38;
		16'h2617: out_word = 8'hCD;
		16'h2618: out_word = 8'hA2;
		16'h2619: out_word = 8'h2D;
		16'h261A: out_word = 8'hED;
		16'h261B: out_word = 8'h43;
		16'h261C: out_word = 8'h76;
		16'h261D: out_word = 8'h5C;
		16'h261E: out_word = 8'h7E;
		16'h261F: out_word = 8'hA7;
		16'h2620: out_word = 8'h28;
		16'h2621: out_word = 8'h03;
		16'h2622: out_word = 8'hD6;
		16'h2623: out_word = 8'h10;
		16'h2624: out_word = 8'h77;
		16'h2625: out_word = 8'h18;
		16'h2626: out_word = 8'h09;
		16'h2627: out_word = 8'hCD;
		16'h2628: out_word = 8'h30;
		16'h2629: out_word = 8'h25;
		16'h262A: out_word = 8'h28;
		16'h262B: out_word = 8'h04;
		16'h262C: out_word = 8'hEF;
		16'h262D: out_word = 8'hA3;
		16'h262E: out_word = 8'h38;
		16'h262F: out_word = 8'h34;
		16'h2630: out_word = 8'hE7;
		16'h2631: out_word = 8'hC3;
		16'h2632: out_word = 8'hC3;
		16'h2633: out_word = 8'h26;
		16'h2634: out_word = 8'h01;
		16'h2635: out_word = 8'h5A;
		16'h2636: out_word = 8'h10;
		16'h2637: out_word = 8'hE7;
		16'h2638: out_word = 8'hFE;
		16'h2639: out_word = 8'h23;
		16'h263A: out_word = 8'hCA;
		16'h263B: out_word = 8'h0D;
		16'h263C: out_word = 8'h27;
		16'h263D: out_word = 8'h21;
		16'h263E: out_word = 8'h3B;
		16'h263F: out_word = 8'h5C;
		16'h2640: out_word = 8'hCB;
		16'h2641: out_word = 8'hB6;
		16'h2642: out_word = 8'hCB;
		16'h2643: out_word = 8'h7E;
		16'h2644: out_word = 8'h28;
		16'h2645: out_word = 8'h1F;
		16'h2646: out_word = 8'hC3;
		16'h2647: out_word = 8'h6C;
		16'h2648: out_word = 8'h3B;
		16'h2649: out_word = 8'h0E;
		16'h264A: out_word = 8'h00;
		16'h264B: out_word = 8'h20;
		16'h264C: out_word = 8'h13;
		16'h264D: out_word = 8'hCD;
		16'h264E: out_word = 8'h1E;
		16'h264F: out_word = 8'h03;
		16'h2650: out_word = 8'h30;
		16'h2651: out_word = 8'h0E;
		16'h2652: out_word = 8'h15;
		16'h2653: out_word = 8'h5F;
		16'h2654: out_word = 8'hCD;
		16'h2655: out_word = 8'h33;
		16'h2656: out_word = 8'h03;
		16'h2657: out_word = 8'hF5;
		16'h2658: out_word = 8'h01;
		16'h2659: out_word = 8'h01;
		16'h265A: out_word = 8'h00;
		16'h265B: out_word = 8'hF7;
		16'h265C: out_word = 8'hF1;
		16'h265D: out_word = 8'h12;
		16'h265E: out_word = 8'h0E;
		16'h265F: out_word = 8'h01;
		16'h2660: out_word = 8'h06;
		16'h2661: out_word = 8'h00;
		16'h2662: out_word = 8'hCD;
		16'h2663: out_word = 8'hB2;
		16'h2664: out_word = 8'h2A;
		16'h2665: out_word = 8'hC3;
		16'h2666: out_word = 8'h12;
		16'h2667: out_word = 8'h27;
		16'h2668: out_word = 8'hCD;
		16'h2669: out_word = 8'h22;
		16'h266A: out_word = 8'h25;
		16'h266B: out_word = 8'hC4;
		16'h266C: out_word = 8'h35;
		16'h266D: out_word = 8'h25;
		16'h266E: out_word = 8'hE7;
		16'h266F: out_word = 8'hC3;
		16'h2670: out_word = 8'hDB;
		16'h2671: out_word = 8'h25;
		16'h2672: out_word = 8'hCD;
		16'h2673: out_word = 8'h22;
		16'h2674: out_word = 8'h25;
		16'h2675: out_word = 8'hC4;
		16'h2676: out_word = 8'h80;
		16'h2677: out_word = 8'h25;
		16'h2678: out_word = 8'hE7;
		16'h2679: out_word = 8'h18;
		16'h267A: out_word = 8'h48;
		16'h267B: out_word = 8'hCD;
		16'h267C: out_word = 8'h22;
		16'h267D: out_word = 8'h25;
		16'h267E: out_word = 8'hC4;
		16'h267F: out_word = 8'hCB;
		16'h2680: out_word = 8'h22;
		16'h2681: out_word = 8'hE7;
		16'h2682: out_word = 8'h18;
		16'h2683: out_word = 8'h3F;
		16'h2684: out_word = 8'hCD;
		16'h2685: out_word = 8'h88;
		16'h2686: out_word = 8'h2C;
		16'h2687: out_word = 8'h30;
		16'h2688: out_word = 8'h56;
		16'h2689: out_word = 8'hFE;
		16'h268A: out_word = 8'h41;
		16'h268B: out_word = 8'h30;
		16'h268C: out_word = 8'h3C;
		16'h268D: out_word = 8'hCD;
		16'h268E: out_word = 8'h30;
		16'h268F: out_word = 8'h25;
		16'h2690: out_word = 8'h20;
		16'h2691: out_word = 8'h23;
		16'h2692: out_word = 8'hCD;
		16'h2693: out_word = 8'h9B;
		16'h2694: out_word = 8'h2C;
		16'h2695: out_word = 8'hDF;
		16'h2696: out_word = 8'h01;
		16'h2697: out_word = 8'h06;
		16'h2698: out_word = 8'h00;
		16'h2699: out_word = 8'hCD;
		16'h269A: out_word = 8'h55;
		16'h269B: out_word = 8'h16;
		16'h269C: out_word = 8'h23;
		16'h269D: out_word = 8'h36;
		16'h269E: out_word = 8'h0E;
		16'h269F: out_word = 8'h23;
		16'h26A0: out_word = 8'hEB;
		16'h26A1: out_word = 8'h2A;
		16'h26A2: out_word = 8'h65;
		16'h26A3: out_word = 8'h5C;
		16'h26A4: out_word = 8'h0E;
		16'h26A5: out_word = 8'h05;
		16'h26A6: out_word = 8'hA7;
		16'h26A7: out_word = 8'hED;
		16'h26A8: out_word = 8'h42;
		16'h26A9: out_word = 8'h22;
		16'h26AA: out_word = 8'h65;
		16'h26AB: out_word = 8'h5C;
		16'h26AC: out_word = 8'hED;
		16'h26AD: out_word = 8'hB0;
		16'h26AE: out_word = 8'hEB;
		16'h26AF: out_word = 8'h2B;
		16'h26B0: out_word = 8'hCD;
		16'h26B1: out_word = 8'h77;
		16'h26B2: out_word = 8'h00;
		16'h26B3: out_word = 8'h18;
		16'h26B4: out_word = 8'h0E;
		16'h26B5: out_word = 8'hDF;
		16'h26B6: out_word = 8'h23;
		16'h26B7: out_word = 8'h7E;
		16'h26B8: out_word = 8'hFE;
		16'h26B9: out_word = 8'h0E;
		16'h26BA: out_word = 8'h20;
		16'h26BB: out_word = 8'hFA;
		16'h26BC: out_word = 8'h23;
		16'h26BD: out_word = 8'hCD;
		16'h26BE: out_word = 8'hB4;
		16'h26BF: out_word = 8'h33;
		16'h26C0: out_word = 8'h22;
		16'h26C1: out_word = 8'h5D;
		16'h26C2: out_word = 8'h5C;
		16'h26C3: out_word = 8'hFD;
		16'h26C4: out_word = 8'hCB;
		16'h26C5: out_word = 8'h01;
		16'h26C6: out_word = 8'hF6;
		16'h26C7: out_word = 8'h18;
		16'h26C8: out_word = 8'h14;
		16'h26C9: out_word = 8'hCD;
		16'h26CA: out_word = 8'hB2;
		16'h26CB: out_word = 8'h28;
		16'h26CC: out_word = 8'hDA;
		16'h26CD: out_word = 8'h2E;
		16'h26CE: out_word = 8'h1C;
		16'h26CF: out_word = 8'hCC;
		16'h26D0: out_word = 8'h96;
		16'h26D1: out_word = 8'h29;
		16'h26D2: out_word = 8'h3A;
		16'h26D3: out_word = 8'h3B;
		16'h26D4: out_word = 8'h5C;
		16'h26D5: out_word = 8'hFE;
		16'h26D6: out_word = 8'hC0;
		16'h26D7: out_word = 8'h38;
		16'h26D8: out_word = 8'h04;
		16'h26D9: out_word = 8'h23;
		16'h26DA: out_word = 8'hCD;
		16'h26DB: out_word = 8'hB4;
		16'h26DC: out_word = 8'h33;
		16'h26DD: out_word = 8'h18;
		16'h26DE: out_word = 8'h33;
		16'h26DF: out_word = 8'h01;
		16'h26E0: out_word = 8'hDB;
		16'h26E1: out_word = 8'h09;
		16'h26E2: out_word = 8'hFE;
		16'h26E3: out_word = 8'h2D;
		16'h26E4: out_word = 8'h28;
		16'h26E5: out_word = 8'h27;
		16'h26E6: out_word = 8'h01;
		16'h26E7: out_word = 8'h18;
		16'h26E8: out_word = 8'h10;
		16'h26E9: out_word = 8'hFE;
		16'h26EA: out_word = 8'hAE;
		16'h26EB: out_word = 8'h28;
		16'h26EC: out_word = 8'h20;
		16'h26ED: out_word = 8'hD6;
		16'h26EE: out_word = 8'hAF;
		16'h26EF: out_word = 8'hDA;
		16'h26F0: out_word = 8'h8A;
		16'h26F1: out_word = 8'h1C;
		16'h26F2: out_word = 8'h01;
		16'h26F3: out_word = 8'hF0;
		16'h26F4: out_word = 8'h04;
		16'h26F5: out_word = 8'hFE;
		16'h26F6: out_word = 8'h14;
		16'h26F7: out_word = 8'h28;
		16'h26F8: out_word = 8'h14;
		16'h26F9: out_word = 8'hD2;
		16'h26FA: out_word = 8'h8A;
		16'h26FB: out_word = 8'h1C;
		16'h26FC: out_word = 8'h06;
		16'h26FD: out_word = 8'h10;
		16'h26FE: out_word = 8'hC6;
		16'h26FF: out_word = 8'hDC;
		16'h2700: out_word = 8'h4F;
		16'h2701: out_word = 8'hFE;
		16'h2702: out_word = 8'hDF;
		16'h2703: out_word = 8'h30;
		16'h2704: out_word = 8'h02;
		16'h2705: out_word = 8'hCB;
		16'h2706: out_word = 8'hB1;
		16'h2707: out_word = 8'hFE;
		16'h2708: out_word = 8'hEE;
		16'h2709: out_word = 8'h38;
		16'h270A: out_word = 8'h02;
		16'h270B: out_word = 8'hCB;
		16'h270C: out_word = 8'hB9;
		16'h270D: out_word = 8'hC5;
		16'h270E: out_word = 8'hE7;
		16'h270F: out_word = 8'hC3;
		16'h2710: out_word = 8'hFF;
		16'h2711: out_word = 8'h24;
		16'h2712: out_word = 8'hDF;
		16'h2713: out_word = 8'hFE;
		16'h2714: out_word = 8'h28;
		16'h2715: out_word = 8'h20;
		16'h2716: out_word = 8'h0C;
		16'h2717: out_word = 8'hFD;
		16'h2718: out_word = 8'hCB;
		16'h2719: out_word = 8'h01;
		16'h271A: out_word = 8'h76;
		16'h271B: out_word = 8'h20;
		16'h271C: out_word = 8'h17;
		16'h271D: out_word = 8'hCD;
		16'h271E: out_word = 8'h52;
		16'h271F: out_word = 8'h2A;
		16'h2720: out_word = 8'hE7;
		16'h2721: out_word = 8'h18;
		16'h2722: out_word = 8'hF0;
		16'h2723: out_word = 8'h06;
		16'h2724: out_word = 8'h00;
		16'h2725: out_word = 8'h4F;
		16'h2726: out_word = 8'h21;
		16'h2727: out_word = 8'h95;
		16'h2728: out_word = 8'h27;
		16'h2729: out_word = 8'hCD;
		16'h272A: out_word = 8'hDC;
		16'h272B: out_word = 8'h16;
		16'h272C: out_word = 8'h30;
		16'h272D: out_word = 8'h06;
		16'h272E: out_word = 8'h4E;
		16'h272F: out_word = 8'h21;
		16'h2730: out_word = 8'hED;
		16'h2731: out_word = 8'h26;
		16'h2732: out_word = 8'h09;
		16'h2733: out_word = 8'h46;
		16'h2734: out_word = 8'hD1;
		16'h2735: out_word = 8'h7A;
		16'h2736: out_word = 8'hB8;
		16'h2737: out_word = 8'h38;
		16'h2738: out_word = 8'h3A;
		16'h2739: out_word = 8'hA7;
		16'h273A: out_word = 8'hCA;
		16'h273B: out_word = 8'h18;
		16'h273C: out_word = 8'h00;
		16'h273D: out_word = 8'hC5;
		16'h273E: out_word = 8'h21;
		16'h273F: out_word = 8'h3B;
		16'h2740: out_word = 8'h5C;
		16'h2741: out_word = 8'h7B;
		16'h2742: out_word = 8'hFE;
		16'h2743: out_word = 8'hED;
		16'h2744: out_word = 8'h20;
		16'h2745: out_word = 8'h06;
		16'h2746: out_word = 8'hCB;
		16'h2747: out_word = 8'h76;
		16'h2748: out_word = 8'h20;
		16'h2749: out_word = 8'h02;
		16'h274A: out_word = 8'h1E;
		16'h274B: out_word = 8'h99;
		16'h274C: out_word = 8'hD5;
		16'h274D: out_word = 8'hCD;
		16'h274E: out_word = 8'h30;
		16'h274F: out_word = 8'h25;
		16'h2750: out_word = 8'h28;
		16'h2751: out_word = 8'h09;
		16'h2752: out_word = 8'h7B;
		16'h2753: out_word = 8'hE6;
		16'h2754: out_word = 8'h3F;
		16'h2755: out_word = 8'h47;
		16'h2756: out_word = 8'hEF;
		16'h2757: out_word = 8'h3B;
		16'h2758: out_word = 8'h38;
		16'h2759: out_word = 8'h18;
		16'h275A: out_word = 8'h09;
		16'h275B: out_word = 8'h7B;
		16'h275C: out_word = 8'hFD;
		16'h275D: out_word = 8'hAE;
		16'h275E: out_word = 8'h01;
		16'h275F: out_word = 8'hE6;
		16'h2760: out_word = 8'h40;
		16'h2761: out_word = 8'hC2;
		16'h2762: out_word = 8'h8A;
		16'h2763: out_word = 8'h1C;
		16'h2764: out_word = 8'hD1;
		16'h2765: out_word = 8'h21;
		16'h2766: out_word = 8'h3B;
		16'h2767: out_word = 8'h5C;
		16'h2768: out_word = 8'hCB;
		16'h2769: out_word = 8'hF6;
		16'h276A: out_word = 8'hCB;
		16'h276B: out_word = 8'h7B;
		16'h276C: out_word = 8'h20;
		16'h276D: out_word = 8'h02;
		16'h276E: out_word = 8'hCB;
		16'h276F: out_word = 8'hB6;
		16'h2770: out_word = 8'hC1;
		16'h2771: out_word = 8'h18;
		16'h2772: out_word = 8'hC1;
		16'h2773: out_word = 8'hD5;
		16'h2774: out_word = 8'h79;
		16'h2775: out_word = 8'hFD;
		16'h2776: out_word = 8'hCB;
		16'h2777: out_word = 8'h01;
		16'h2778: out_word = 8'h76;
		16'h2779: out_word = 8'h20;
		16'h277A: out_word = 8'h15;
		16'h277B: out_word = 8'hE6;
		16'h277C: out_word = 8'h3F;
		16'h277D: out_word = 8'hC6;
		16'h277E: out_word = 8'h08;
		16'h277F: out_word = 8'h4F;
		16'h2780: out_word = 8'hFE;
		16'h2781: out_word = 8'h10;
		16'h2782: out_word = 8'h20;
		16'h2783: out_word = 8'h04;
		16'h2784: out_word = 8'hCB;
		16'h2785: out_word = 8'hF1;
		16'h2786: out_word = 8'h18;
		16'h2787: out_word = 8'h08;
		16'h2788: out_word = 8'h38;
		16'h2789: out_word = 8'hD7;
		16'h278A: out_word = 8'hFE;
		16'h278B: out_word = 8'h17;
		16'h278C: out_word = 8'h28;
		16'h278D: out_word = 8'h02;
		16'h278E: out_word = 8'hCB;
		16'h278F: out_word = 8'hF9;
		16'h2790: out_word = 8'hC5;
		16'h2791: out_word = 8'hE7;
		16'h2792: out_word = 8'hC3;
		16'h2793: out_word = 8'hFF;
		16'h2794: out_word = 8'h24;
		16'h2795: out_word = 8'h2B;
		16'h2796: out_word = 8'hCF;
		16'h2797: out_word = 8'h2D;
		16'h2798: out_word = 8'hC3;
		16'h2799: out_word = 8'h2A;
		16'h279A: out_word = 8'hC4;
		16'h279B: out_word = 8'h2F;
		16'h279C: out_word = 8'hC5;
		16'h279D: out_word = 8'h5E;
		16'h279E: out_word = 8'hC6;
		16'h279F: out_word = 8'h3D;
		16'h27A0: out_word = 8'hCE;
		16'h27A1: out_word = 8'h3E;
		16'h27A2: out_word = 8'hCC;
		16'h27A3: out_word = 8'h3C;
		16'h27A4: out_word = 8'hCD;
		16'h27A5: out_word = 8'hC7;
		16'h27A6: out_word = 8'hC9;
		16'h27A7: out_word = 8'hC8;
		16'h27A8: out_word = 8'hCA;
		16'h27A9: out_word = 8'hC9;
		16'h27AA: out_word = 8'hCB;
		16'h27AB: out_word = 8'hC5;
		16'h27AC: out_word = 8'hC7;
		16'h27AD: out_word = 8'hC6;
		16'h27AE: out_word = 8'hC8;
		16'h27AF: out_word = 8'h00;
		16'h27B0: out_word = 8'h06;
		16'h27B1: out_word = 8'h08;
		16'h27B2: out_word = 8'h08;
		16'h27B3: out_word = 8'h0A;
		16'h27B4: out_word = 8'h02;
		16'h27B5: out_word = 8'h03;
		16'h27B6: out_word = 8'h05;
		16'h27B7: out_word = 8'h05;
		16'h27B8: out_word = 8'h05;
		16'h27B9: out_word = 8'h05;
		16'h27BA: out_word = 8'h05;
		16'h27BB: out_word = 8'h05;
		16'h27BC: out_word = 8'h06;
		16'h27BD: out_word = 8'hCD;
		16'h27BE: out_word = 8'h30;
		16'h27BF: out_word = 8'h25;
		16'h27C0: out_word = 8'h20;
		16'h27C1: out_word = 8'h35;
		16'h27C2: out_word = 8'hE7;
		16'h27C3: out_word = 8'hCD;
		16'h27C4: out_word = 8'h8D;
		16'h27C5: out_word = 8'h2C;
		16'h27C6: out_word = 8'hD2;
		16'h27C7: out_word = 8'h8A;
		16'h27C8: out_word = 8'h1C;
		16'h27C9: out_word = 8'hE7;
		16'h27CA: out_word = 8'hFE;
		16'h27CB: out_word = 8'h24;
		16'h27CC: out_word = 8'hF5;
		16'h27CD: out_word = 8'h20;
		16'h27CE: out_word = 8'h01;
		16'h27CF: out_word = 8'hE7;
		16'h27D0: out_word = 8'hFE;
		16'h27D1: out_word = 8'h28;
		16'h27D2: out_word = 8'h20;
		16'h27D3: out_word = 8'h12;
		16'h27D4: out_word = 8'hE7;
		16'h27D5: out_word = 8'hFE;
		16'h27D6: out_word = 8'h29;
		16'h27D7: out_word = 8'h28;
		16'h27D8: out_word = 8'h10;
		16'h27D9: out_word = 8'hCD;
		16'h27DA: out_word = 8'hFB;
		16'h27DB: out_word = 8'h24;
		16'h27DC: out_word = 8'hDF;
		16'h27DD: out_word = 8'hFE;
		16'h27DE: out_word = 8'h2C;
		16'h27DF: out_word = 8'h20;
		16'h27E0: out_word = 8'h03;
		16'h27E1: out_word = 8'hE7;
		16'h27E2: out_word = 8'h18;
		16'h27E3: out_word = 8'hF5;
		16'h27E4: out_word = 8'hFE;
		16'h27E5: out_word = 8'h29;
		16'h27E6: out_word = 8'hC2;
		16'h27E7: out_word = 8'h8A;
		16'h27E8: out_word = 8'h1C;
		16'h27E9: out_word = 8'hE7;
		16'h27EA: out_word = 8'h21;
		16'h27EB: out_word = 8'h3B;
		16'h27EC: out_word = 8'h5C;
		16'h27ED: out_word = 8'hCB;
		16'h27EE: out_word = 8'hB6;
		16'h27EF: out_word = 8'hF1;
		16'h27F0: out_word = 8'h28;
		16'h27F1: out_word = 8'h02;
		16'h27F2: out_word = 8'hCB;
		16'h27F3: out_word = 8'hF6;
		16'h27F4: out_word = 8'hC3;
		16'h27F5: out_word = 8'h12;
		16'h27F6: out_word = 8'h27;
		16'h27F7: out_word = 8'hE7;
		16'h27F8: out_word = 8'hE6;
		16'h27F9: out_word = 8'hDF;
		16'h27FA: out_word = 8'h47;
		16'h27FB: out_word = 8'hE7;
		16'h27FC: out_word = 8'hD6;
		16'h27FD: out_word = 8'h24;
		16'h27FE: out_word = 8'h4F;
		16'h27FF: out_word = 8'h20;
		16'h2800: out_word = 8'h01;
		16'h2801: out_word = 8'hE7;
		16'h2802: out_word = 8'hE7;
		16'h2803: out_word = 8'hE5;
		16'h2804: out_word = 8'h2A;
		16'h2805: out_word = 8'h53;
		16'h2806: out_word = 8'h5C;
		16'h2807: out_word = 8'h2B;
		16'h2808: out_word = 8'h11;
		16'h2809: out_word = 8'hCE;
		16'h280A: out_word = 8'h00;
		16'h280B: out_word = 8'hC5;
		16'h280C: out_word = 8'hCD;
		16'h280D: out_word = 8'h86;
		16'h280E: out_word = 8'h1D;
		16'h280F: out_word = 8'hC1;
		16'h2810: out_word = 8'h30;
		16'h2811: out_word = 8'h02;
		16'h2812: out_word = 8'hCF;
		16'h2813: out_word = 8'h18;
		16'h2814: out_word = 8'hE5;
		16'h2815: out_word = 8'hCD;
		16'h2816: out_word = 8'hAB;
		16'h2817: out_word = 8'h28;
		16'h2818: out_word = 8'hE6;
		16'h2819: out_word = 8'hDF;
		16'h281A: out_word = 8'hB8;
		16'h281B: out_word = 8'h20;
		16'h281C: out_word = 8'h08;
		16'h281D: out_word = 8'hCD;
		16'h281E: out_word = 8'hAB;
		16'h281F: out_word = 8'h28;
		16'h2820: out_word = 8'hD6;
		16'h2821: out_word = 8'h24;
		16'h2822: out_word = 8'hB9;
		16'h2823: out_word = 8'h28;
		16'h2824: out_word = 8'h0C;
		16'h2825: out_word = 8'hE1;
		16'h2826: out_word = 8'h2B;
		16'h2827: out_word = 8'h11;
		16'h2828: out_word = 8'h00;
		16'h2829: out_word = 8'h02;
		16'h282A: out_word = 8'hC5;
		16'h282B: out_word = 8'hCD;
		16'h282C: out_word = 8'h8B;
		16'h282D: out_word = 8'h19;
		16'h282E: out_word = 8'hC1;
		16'h282F: out_word = 8'h18;
		16'h2830: out_word = 8'hD7;
		16'h2831: out_word = 8'hA7;
		16'h2832: out_word = 8'hCC;
		16'h2833: out_word = 8'hAB;
		16'h2834: out_word = 8'h28;
		16'h2835: out_word = 8'hD1;
		16'h2836: out_word = 8'hD1;
		16'h2837: out_word = 8'hED;
		16'h2838: out_word = 8'h53;
		16'h2839: out_word = 8'h5D;
		16'h283A: out_word = 8'h5C;
		16'h283B: out_word = 8'hCD;
		16'h283C: out_word = 8'hAB;
		16'h283D: out_word = 8'h28;
		16'h283E: out_word = 8'hE5;
		16'h283F: out_word = 8'hFE;
		16'h2840: out_word = 8'h29;
		16'h2841: out_word = 8'h28;
		16'h2842: out_word = 8'h42;
		16'h2843: out_word = 8'h23;
		16'h2844: out_word = 8'h7E;
		16'h2845: out_word = 8'hFE;
		16'h2846: out_word = 8'h0E;
		16'h2847: out_word = 8'h16;
		16'h2848: out_word = 8'h40;
		16'h2849: out_word = 8'h28;
		16'h284A: out_word = 8'h07;
		16'h284B: out_word = 8'h2B;
		16'h284C: out_word = 8'hCD;
		16'h284D: out_word = 8'hAB;
		16'h284E: out_word = 8'h28;
		16'h284F: out_word = 8'h23;
		16'h2850: out_word = 8'h16;
		16'h2851: out_word = 8'h00;
		16'h2852: out_word = 8'h23;
		16'h2853: out_word = 8'hE5;
		16'h2854: out_word = 8'hD5;
		16'h2855: out_word = 8'hCD;
		16'h2856: out_word = 8'hFB;
		16'h2857: out_word = 8'h24;
		16'h2858: out_word = 8'hF1;
		16'h2859: out_word = 8'hFD;
		16'h285A: out_word = 8'hAE;
		16'h285B: out_word = 8'h01;
		16'h285C: out_word = 8'hE6;
		16'h285D: out_word = 8'h40;
		16'h285E: out_word = 8'h20;
		16'h285F: out_word = 8'h2B;
		16'h2860: out_word = 8'hE1;
		16'h2861: out_word = 8'hEB;
		16'h2862: out_word = 8'h2A;
		16'h2863: out_word = 8'h65;
		16'h2864: out_word = 8'h5C;
		16'h2865: out_word = 8'h01;
		16'h2866: out_word = 8'h05;
		16'h2867: out_word = 8'h00;
		16'h2868: out_word = 8'hED;
		16'h2869: out_word = 8'h42;
		16'h286A: out_word = 8'h22;
		16'h286B: out_word = 8'h65;
		16'h286C: out_word = 8'h5C;
		16'h286D: out_word = 8'hED;
		16'h286E: out_word = 8'hB0;
		16'h286F: out_word = 8'hEB;
		16'h2870: out_word = 8'h2B;
		16'h2871: out_word = 8'hCD;
		16'h2872: out_word = 8'hAB;
		16'h2873: out_word = 8'h28;
		16'h2874: out_word = 8'hFE;
		16'h2875: out_word = 8'h29;
		16'h2876: out_word = 8'h28;
		16'h2877: out_word = 8'h0D;
		16'h2878: out_word = 8'hE5;
		16'h2879: out_word = 8'hDF;
		16'h287A: out_word = 8'hFE;
		16'h287B: out_word = 8'h2C;
		16'h287C: out_word = 8'h20;
		16'h287D: out_word = 8'h0D;
		16'h287E: out_word = 8'hE7;
		16'h287F: out_word = 8'hE1;
		16'h2880: out_word = 8'hCD;
		16'h2881: out_word = 8'hAB;
		16'h2882: out_word = 8'h28;
		16'h2883: out_word = 8'h18;
		16'h2884: out_word = 8'hBE;
		16'h2885: out_word = 8'hE5;
		16'h2886: out_word = 8'hDF;
		16'h2887: out_word = 8'hFE;
		16'h2888: out_word = 8'h29;
		16'h2889: out_word = 8'h28;
		16'h288A: out_word = 8'h02;
		16'h288B: out_word = 8'hCF;
		16'h288C: out_word = 8'h19;
		16'h288D: out_word = 8'hD1;
		16'h288E: out_word = 8'hEB;
		16'h288F: out_word = 8'h22;
		16'h2890: out_word = 8'h5D;
		16'h2891: out_word = 8'h5C;
		16'h2892: out_word = 8'h2A;
		16'h2893: out_word = 8'h0B;
		16'h2894: out_word = 8'h5C;
		16'h2895: out_word = 8'hE3;
		16'h2896: out_word = 8'h22;
		16'h2897: out_word = 8'h0B;
		16'h2898: out_word = 8'h5C;
		16'h2899: out_word = 8'hD5;
		16'h289A: out_word = 8'hE7;
		16'h289B: out_word = 8'hE7;
		16'h289C: out_word = 8'hCD;
		16'h289D: out_word = 8'hFB;
		16'h289E: out_word = 8'h24;
		16'h289F: out_word = 8'hE1;
		16'h28A0: out_word = 8'h22;
		16'h28A1: out_word = 8'h5D;
		16'h28A2: out_word = 8'h5C;
		16'h28A3: out_word = 8'hE1;
		16'h28A4: out_word = 8'h22;
		16'h28A5: out_word = 8'h0B;
		16'h28A6: out_word = 8'h5C;
		16'h28A7: out_word = 8'hE7;
		16'h28A8: out_word = 8'hC3;
		16'h28A9: out_word = 8'h12;
		16'h28AA: out_word = 8'h27;
		16'h28AB: out_word = 8'h23;
		16'h28AC: out_word = 8'h7E;
		16'h28AD: out_word = 8'hFE;
		16'h28AE: out_word = 8'h21;
		16'h28AF: out_word = 8'h38;
		16'h28B0: out_word = 8'hFA;
		16'h28B1: out_word = 8'hC9;
		16'h28B2: out_word = 8'hFD;
		16'h28B3: out_word = 8'hCB;
		16'h28B4: out_word = 8'h01;
		16'h28B5: out_word = 8'hF6;
		16'h28B6: out_word = 8'hDF;
		16'h28B7: out_word = 8'hCD;
		16'h28B8: out_word = 8'h8D;
		16'h28B9: out_word = 8'h2C;
		16'h28BA: out_word = 8'hD2;
		16'h28BB: out_word = 8'h8A;
		16'h28BC: out_word = 8'h1C;
		16'h28BD: out_word = 8'hE5;
		16'h28BE: out_word = 8'hE6;
		16'h28BF: out_word = 8'h1F;
		16'h28C0: out_word = 8'h4F;
		16'h28C1: out_word = 8'hE7;
		16'h28C2: out_word = 8'hE5;
		16'h28C3: out_word = 8'hFE;
		16'h28C4: out_word = 8'h28;
		16'h28C5: out_word = 8'h28;
		16'h28C6: out_word = 8'h28;
		16'h28C7: out_word = 8'hCB;
		16'h28C8: out_word = 8'hF1;
		16'h28C9: out_word = 8'hFE;
		16'h28CA: out_word = 8'h24;
		16'h28CB: out_word = 8'h28;
		16'h28CC: out_word = 8'h11;
		16'h28CD: out_word = 8'hCB;
		16'h28CE: out_word = 8'hE9;
		16'h28CF: out_word = 8'hCD;
		16'h28D0: out_word = 8'h88;
		16'h28D1: out_word = 8'h2C;
		16'h28D2: out_word = 8'h30;
		16'h28D3: out_word = 8'h0F;
		16'h28D4: out_word = 8'hCD;
		16'h28D5: out_word = 8'h88;
		16'h28D6: out_word = 8'h2C;
		16'h28D7: out_word = 8'h30;
		16'h28D8: out_word = 8'h16;
		16'h28D9: out_word = 8'hCB;
		16'h28DA: out_word = 8'hB1;
		16'h28DB: out_word = 8'hE7;
		16'h28DC: out_word = 8'h18;
		16'h28DD: out_word = 8'hF6;
		16'h28DE: out_word = 8'hE7;
		16'h28DF: out_word = 8'hFD;
		16'h28E0: out_word = 8'hCB;
		16'h28E1: out_word = 8'h01;
		16'h28E2: out_word = 8'hB6;
		16'h28E3: out_word = 8'h3A;
		16'h28E4: out_word = 8'h0C;
		16'h28E5: out_word = 8'h5C;
		16'h28E6: out_word = 8'hA7;
		16'h28E7: out_word = 8'h28;
		16'h28E8: out_word = 8'h06;
		16'h28E9: out_word = 8'hCD;
		16'h28EA: out_word = 8'h30;
		16'h28EB: out_word = 8'h25;
		16'h28EC: out_word = 8'hC2;
		16'h28ED: out_word = 8'h51;
		16'h28EE: out_word = 8'h29;
		16'h28EF: out_word = 8'h41;
		16'h28F0: out_word = 8'hCD;
		16'h28F1: out_word = 8'h30;
		16'h28F2: out_word = 8'h25;
		16'h28F3: out_word = 8'h20;
		16'h28F4: out_word = 8'h08;
		16'h28F5: out_word = 8'h79;
		16'h28F6: out_word = 8'hE6;
		16'h28F7: out_word = 8'hE0;
		16'h28F8: out_word = 8'hCB;
		16'h28F9: out_word = 8'hFF;
		16'h28FA: out_word = 8'h4F;
		16'h28FB: out_word = 8'h18;
		16'h28FC: out_word = 8'h37;
		16'h28FD: out_word = 8'h2A;
		16'h28FE: out_word = 8'h4B;
		16'h28FF: out_word = 8'h5C;
		16'h2900: out_word = 8'h7E;
		16'h2901: out_word = 8'hE6;
		16'h2902: out_word = 8'h7F;
		16'h2903: out_word = 8'h28;
		16'h2904: out_word = 8'h2D;
		16'h2905: out_word = 8'hB9;
		16'h2906: out_word = 8'h20;
		16'h2907: out_word = 8'h22;
		16'h2908: out_word = 8'h17;
		16'h2909: out_word = 8'h87;
		16'h290A: out_word = 8'hF2;
		16'h290B: out_word = 8'h3F;
		16'h290C: out_word = 8'h29;
		16'h290D: out_word = 8'h38;
		16'h290E: out_word = 8'h30;
		16'h290F: out_word = 8'hD1;
		16'h2910: out_word = 8'hD5;
		16'h2911: out_word = 8'hE5;
		16'h2912: out_word = 8'h23;
		16'h2913: out_word = 8'h1A;
		16'h2914: out_word = 8'h13;
		16'h2915: out_word = 8'hFE;
		16'h2916: out_word = 8'h20;
		16'h2917: out_word = 8'h28;
		16'h2918: out_word = 8'hFA;
		16'h2919: out_word = 8'hF6;
		16'h291A: out_word = 8'h20;
		16'h291B: out_word = 8'hBE;
		16'h291C: out_word = 8'h28;
		16'h291D: out_word = 8'hF4;
		16'h291E: out_word = 8'hF6;
		16'h291F: out_word = 8'h80;
		16'h2920: out_word = 8'hBE;
		16'h2921: out_word = 8'h20;
		16'h2922: out_word = 8'h06;
		16'h2923: out_word = 8'h1A;
		16'h2924: out_word = 8'hCD;
		16'h2925: out_word = 8'h88;
		16'h2926: out_word = 8'h2C;
		16'h2927: out_word = 8'h30;
		16'h2928: out_word = 8'h15;
		16'h2929: out_word = 8'hE1;
		16'h292A: out_word = 8'hC5;
		16'h292B: out_word = 8'hCD;
		16'h292C: out_word = 8'hB8;
		16'h292D: out_word = 8'h19;
		16'h292E: out_word = 8'hEB;
		16'h292F: out_word = 8'hC1;
		16'h2930: out_word = 8'h18;
		16'h2931: out_word = 8'hCE;
		16'h2932: out_word = 8'hCB;
		16'h2933: out_word = 8'hF8;
		16'h2934: out_word = 8'hD1;
		16'h2935: out_word = 8'hDF;
		16'h2936: out_word = 8'hFE;
		16'h2937: out_word = 8'h28;
		16'h2938: out_word = 8'h28;
		16'h2939: out_word = 8'h09;
		16'h293A: out_word = 8'hCB;
		16'h293B: out_word = 8'hE8;
		16'h293C: out_word = 8'h18;
		16'h293D: out_word = 8'h0D;
		16'h293E: out_word = 8'hD1;
		16'h293F: out_word = 8'hD1;
		16'h2940: out_word = 8'hD1;
		16'h2941: out_word = 8'hE5;
		16'h2942: out_word = 8'hDF;
		16'h2943: out_word = 8'hCD;
		16'h2944: out_word = 8'h88;
		16'h2945: out_word = 8'h2C;
		16'h2946: out_word = 8'h30;
		16'h2947: out_word = 8'h03;
		16'h2948: out_word = 8'hE7;
		16'h2949: out_word = 8'h18;
		16'h294A: out_word = 8'hF8;
		16'h294B: out_word = 8'hE1;
		16'h294C: out_word = 8'hCB;
		16'h294D: out_word = 8'h10;
		16'h294E: out_word = 8'hCB;
		16'h294F: out_word = 8'h70;
		16'h2950: out_word = 8'hC9;
		16'h2951: out_word = 8'h2A;
		16'h2952: out_word = 8'h0B;
		16'h2953: out_word = 8'h5C;
		16'h2954: out_word = 8'h7E;
		16'h2955: out_word = 8'hFE;
		16'h2956: out_word = 8'h29;
		16'h2957: out_word = 8'hCA;
		16'h2958: out_word = 8'hEF;
		16'h2959: out_word = 8'h28;
		16'h295A: out_word = 8'h7E;
		16'h295B: out_word = 8'hF6;
		16'h295C: out_word = 8'h60;
		16'h295D: out_word = 8'h47;
		16'h295E: out_word = 8'h23;
		16'h295F: out_word = 8'h7E;
		16'h2960: out_word = 8'hFE;
		16'h2961: out_word = 8'h0E;
		16'h2962: out_word = 8'h28;
		16'h2963: out_word = 8'h07;
		16'h2964: out_word = 8'h2B;
		16'h2965: out_word = 8'hCD;
		16'h2966: out_word = 8'hAB;
		16'h2967: out_word = 8'h28;
		16'h2968: out_word = 8'h23;
		16'h2969: out_word = 8'hCB;
		16'h296A: out_word = 8'hA8;
		16'h296B: out_word = 8'h78;
		16'h296C: out_word = 8'hB9;
		16'h296D: out_word = 8'h28;
		16'h296E: out_word = 8'h12;
		16'h296F: out_word = 8'h23;
		16'h2970: out_word = 8'h23;
		16'h2971: out_word = 8'h23;
		16'h2972: out_word = 8'h23;
		16'h2973: out_word = 8'h23;
		16'h2974: out_word = 8'hCD;
		16'h2975: out_word = 8'hAB;
		16'h2976: out_word = 8'h28;
		16'h2977: out_word = 8'hFE;
		16'h2978: out_word = 8'h29;
		16'h2979: out_word = 8'hCA;
		16'h297A: out_word = 8'hEF;
		16'h297B: out_word = 8'h28;
		16'h297C: out_word = 8'hCD;
		16'h297D: out_word = 8'hAB;
		16'h297E: out_word = 8'h28;
		16'h297F: out_word = 8'h18;
		16'h2980: out_word = 8'hD9;
		16'h2981: out_word = 8'hCB;
		16'h2982: out_word = 8'h69;
		16'h2983: out_word = 8'h20;
		16'h2984: out_word = 8'h0C;
		16'h2985: out_word = 8'h23;
		16'h2986: out_word = 8'hED;
		16'h2987: out_word = 8'h5B;
		16'h2988: out_word = 8'h65;
		16'h2989: out_word = 8'h5C;
		16'h298A: out_word = 8'hCD;
		16'h298B: out_word = 8'hC0;
		16'h298C: out_word = 8'h33;
		16'h298D: out_word = 8'hEB;
		16'h298E: out_word = 8'h22;
		16'h298F: out_word = 8'h65;
		16'h2990: out_word = 8'h5C;
		16'h2991: out_word = 8'hD1;
		16'h2992: out_word = 8'hD1;
		16'h2993: out_word = 8'hAF;
		16'h2994: out_word = 8'h3C;
		16'h2995: out_word = 8'hC9;
		16'h2996: out_word = 8'hAF;
		16'h2997: out_word = 8'h47;
		16'h2998: out_word = 8'hCB;
		16'h2999: out_word = 8'h79;
		16'h299A: out_word = 8'h20;
		16'h299B: out_word = 8'h4B;
		16'h299C: out_word = 8'hCB;
		16'h299D: out_word = 8'h7E;
		16'h299E: out_word = 8'h20;
		16'h299F: out_word = 8'h0E;
		16'h29A0: out_word = 8'h3C;
		16'h29A1: out_word = 8'h23;
		16'h29A2: out_word = 8'h4E;
		16'h29A3: out_word = 8'h23;
		16'h29A4: out_word = 8'h46;
		16'h29A5: out_word = 8'h23;
		16'h29A6: out_word = 8'hEB;
		16'h29A7: out_word = 8'hCD;
		16'h29A8: out_word = 8'hB2;
		16'h29A9: out_word = 8'h2A;
		16'h29AA: out_word = 8'hDF;
		16'h29AB: out_word = 8'hC3;
		16'h29AC: out_word = 8'h49;
		16'h29AD: out_word = 8'h2A;
		16'h29AE: out_word = 8'h23;
		16'h29AF: out_word = 8'h23;
		16'h29B0: out_word = 8'h23;
		16'h29B1: out_word = 8'h46;
		16'h29B2: out_word = 8'hCB;
		16'h29B3: out_word = 8'h71;
		16'h29B4: out_word = 8'h28;
		16'h29B5: out_word = 8'h0A;
		16'h29B6: out_word = 8'h05;
		16'h29B7: out_word = 8'h28;
		16'h29B8: out_word = 8'hE8;
		16'h29B9: out_word = 8'hEB;
		16'h29BA: out_word = 8'hDF;
		16'h29BB: out_word = 8'hFE;
		16'h29BC: out_word = 8'h28;
		16'h29BD: out_word = 8'h20;
		16'h29BE: out_word = 8'h61;
		16'h29BF: out_word = 8'hEB;
		16'h29C0: out_word = 8'hEB;
		16'h29C1: out_word = 8'h18;
		16'h29C2: out_word = 8'h24;
		16'h29C3: out_word = 8'hE5;
		16'h29C4: out_word = 8'hDF;
		16'h29C5: out_word = 8'hE1;
		16'h29C6: out_word = 8'hFE;
		16'h29C7: out_word = 8'h2C;
		16'h29C8: out_word = 8'h28;
		16'h29C9: out_word = 8'h20;
		16'h29CA: out_word = 8'hCB;
		16'h29CB: out_word = 8'h79;
		16'h29CC: out_word = 8'h28;
		16'h29CD: out_word = 8'h52;
		16'h29CE: out_word = 8'hCB;
		16'h29CF: out_word = 8'h71;
		16'h29D0: out_word = 8'h20;
		16'h29D1: out_word = 8'h06;
		16'h29D2: out_word = 8'hFE;
		16'h29D3: out_word = 8'h29;
		16'h29D4: out_word = 8'h20;
		16'h29D5: out_word = 8'h3C;
		16'h29D6: out_word = 8'hE7;
		16'h29D7: out_word = 8'hC9;
		16'h29D8: out_word = 8'hFE;
		16'h29D9: out_word = 8'h29;
		16'h29DA: out_word = 8'h28;
		16'h29DB: out_word = 8'h6C;
		16'h29DC: out_word = 8'hFE;
		16'h29DD: out_word = 8'hCC;
		16'h29DE: out_word = 8'h20;
		16'h29DF: out_word = 8'h32;
		16'h29E0: out_word = 8'hDF;
		16'h29E1: out_word = 8'h2B;
		16'h29E2: out_word = 8'h22;
		16'h29E3: out_word = 8'h5D;
		16'h29E4: out_word = 8'h5C;
		16'h29E5: out_word = 8'h18;
		16'h29E6: out_word = 8'h5E;
		16'h29E7: out_word = 8'h21;
		16'h29E8: out_word = 8'h00;
		16'h29E9: out_word = 8'h00;
		16'h29EA: out_word = 8'hE5;
		16'h29EB: out_word = 8'hE7;
		16'h29EC: out_word = 8'hE1;
		16'h29ED: out_word = 8'h79;
		16'h29EE: out_word = 8'hFE;
		16'h29EF: out_word = 8'hC0;
		16'h29F0: out_word = 8'h20;
		16'h29F1: out_word = 8'h09;
		16'h29F2: out_word = 8'hDF;
		16'h29F3: out_word = 8'hFE;
		16'h29F4: out_word = 8'h29;
		16'h29F5: out_word = 8'h28;
		16'h29F6: out_word = 8'h51;
		16'h29F7: out_word = 8'hFE;
		16'h29F8: out_word = 8'hCC;
		16'h29F9: out_word = 8'h28;
		16'h29FA: out_word = 8'hE5;
		16'h29FB: out_word = 8'hC5;
		16'h29FC: out_word = 8'hE5;
		16'h29FD: out_word = 8'hCD;
		16'h29FE: out_word = 8'hEE;
		16'h29FF: out_word = 8'h2A;
		16'h2A00: out_word = 8'hE3;
		16'h2A01: out_word = 8'hEB;
		16'h2A02: out_word = 8'hCD;
		16'h2A03: out_word = 8'hCC;
		16'h2A04: out_word = 8'h2A;
		16'h2A05: out_word = 8'h38;
		16'h2A06: out_word = 8'h19;
		16'h2A07: out_word = 8'h0B;
		16'h2A08: out_word = 8'hCD;
		16'h2A09: out_word = 8'hF4;
		16'h2A0A: out_word = 8'h2A;
		16'h2A0B: out_word = 8'h09;
		16'h2A0C: out_word = 8'hD1;
		16'h2A0D: out_word = 8'hC1;
		16'h2A0E: out_word = 8'h10;
		16'h2A0F: out_word = 8'hB3;
		16'h2A10: out_word = 8'hCB;
		16'h2A11: out_word = 8'h79;
		16'h2A12: out_word = 8'h20;
		16'h2A13: out_word = 8'h66;
		16'h2A14: out_word = 8'hE5;
		16'h2A15: out_word = 8'hCB;
		16'h2A16: out_word = 8'h71;
		16'h2A17: out_word = 8'h20;
		16'h2A18: out_word = 8'h13;
		16'h2A19: out_word = 8'h42;
		16'h2A1A: out_word = 8'h4B;
		16'h2A1B: out_word = 8'hDF;
		16'h2A1C: out_word = 8'hFE;
		16'h2A1D: out_word = 8'h29;
		16'h2A1E: out_word = 8'h28;
		16'h2A1F: out_word = 8'h02;
		16'h2A20: out_word = 8'hCF;
		16'h2A21: out_word = 8'h02;
		16'h2A22: out_word = 8'hE7;
		16'h2A23: out_word = 8'hE1;
		16'h2A24: out_word = 8'h11;
		16'h2A25: out_word = 8'h05;
		16'h2A26: out_word = 8'h00;
		16'h2A27: out_word = 8'hCD;
		16'h2A28: out_word = 8'hF4;
		16'h2A29: out_word = 8'h2A;
		16'h2A2A: out_word = 8'h09;
		16'h2A2B: out_word = 8'hC9;
		16'h2A2C: out_word = 8'hCD;
		16'h2A2D: out_word = 8'hEE;
		16'h2A2E: out_word = 8'h2A;
		16'h2A2F: out_word = 8'hE3;
		16'h2A30: out_word = 8'hCD;
		16'h2A31: out_word = 8'hF4;
		16'h2A32: out_word = 8'h2A;
		16'h2A33: out_word = 8'hC1;
		16'h2A34: out_word = 8'h09;
		16'h2A35: out_word = 8'h23;
		16'h2A36: out_word = 8'h42;
		16'h2A37: out_word = 8'h4B;
		16'h2A38: out_word = 8'hEB;
		16'h2A39: out_word = 8'hCD;
		16'h2A3A: out_word = 8'hB1;
		16'h2A3B: out_word = 8'h2A;
		16'h2A3C: out_word = 8'hDF;
		16'h2A3D: out_word = 8'hFE;
		16'h2A3E: out_word = 8'h29;
		16'h2A3F: out_word = 8'h28;
		16'h2A40: out_word = 8'h07;
		16'h2A41: out_word = 8'hFE;
		16'h2A42: out_word = 8'h2C;
		16'h2A43: out_word = 8'h20;
		16'h2A44: out_word = 8'hDB;
		16'h2A45: out_word = 8'hCD;
		16'h2A46: out_word = 8'h52;
		16'h2A47: out_word = 8'h2A;
		16'h2A48: out_word = 8'hE7;
		16'h2A49: out_word = 8'hFE;
		16'h2A4A: out_word = 8'h28;
		16'h2A4B: out_word = 8'h28;
		16'h2A4C: out_word = 8'hF8;
		16'h2A4D: out_word = 8'hFD;
		16'h2A4E: out_word = 8'hCB;
		16'h2A4F: out_word = 8'h01;
		16'h2A50: out_word = 8'hB6;
		16'h2A51: out_word = 8'hC9;
		16'h2A52: out_word = 8'hCD;
		16'h2A53: out_word = 8'h30;
		16'h2A54: out_word = 8'h25;
		16'h2A55: out_word = 8'hC4;
		16'h2A56: out_word = 8'hF1;
		16'h2A57: out_word = 8'h2B;
		16'h2A58: out_word = 8'hE7;
		16'h2A59: out_word = 8'hFE;
		16'h2A5A: out_word = 8'h29;
		16'h2A5B: out_word = 8'h28;
		16'h2A5C: out_word = 8'h50;
		16'h2A5D: out_word = 8'hD5;
		16'h2A5E: out_word = 8'hAF;
		16'h2A5F: out_word = 8'hF5;
		16'h2A60: out_word = 8'hC5;
		16'h2A61: out_word = 8'h11;
		16'h2A62: out_word = 8'h01;
		16'h2A63: out_word = 8'h00;
		16'h2A64: out_word = 8'hDF;
		16'h2A65: out_word = 8'hE1;
		16'h2A66: out_word = 8'hFE;
		16'h2A67: out_word = 8'hCC;
		16'h2A68: out_word = 8'h28;
		16'h2A69: out_word = 8'h17;
		16'h2A6A: out_word = 8'hF1;
		16'h2A6B: out_word = 8'hCD;
		16'h2A6C: out_word = 8'hCD;
		16'h2A6D: out_word = 8'h2A;
		16'h2A6E: out_word = 8'hF5;
		16'h2A6F: out_word = 8'h50;
		16'h2A70: out_word = 8'h59;
		16'h2A71: out_word = 8'hE5;
		16'h2A72: out_word = 8'hDF;
		16'h2A73: out_word = 8'hE1;
		16'h2A74: out_word = 8'hFE;
		16'h2A75: out_word = 8'hCC;
		16'h2A76: out_word = 8'h28;
		16'h2A77: out_word = 8'h09;
		16'h2A78: out_word = 8'hFE;
		16'h2A79: out_word = 8'h29;
		16'h2A7A: out_word = 8'hC2;
		16'h2A7B: out_word = 8'h8A;
		16'h2A7C: out_word = 8'h1C;
		16'h2A7D: out_word = 8'h62;
		16'h2A7E: out_word = 8'h6B;
		16'h2A7F: out_word = 8'h18;
		16'h2A80: out_word = 8'h13;
		16'h2A81: out_word = 8'hE5;
		16'h2A82: out_word = 8'hE7;
		16'h2A83: out_word = 8'hE1;
		16'h2A84: out_word = 8'hFE;
		16'h2A85: out_word = 8'h29;
		16'h2A86: out_word = 8'h28;
		16'h2A87: out_word = 8'h0C;
		16'h2A88: out_word = 8'hF1;
		16'h2A89: out_word = 8'hCD;
		16'h2A8A: out_word = 8'hCD;
		16'h2A8B: out_word = 8'h2A;
		16'h2A8C: out_word = 8'hF5;
		16'h2A8D: out_word = 8'hDF;
		16'h2A8E: out_word = 8'h60;
		16'h2A8F: out_word = 8'h69;
		16'h2A90: out_word = 8'hFE;
		16'h2A91: out_word = 8'h29;
		16'h2A92: out_word = 8'h20;
		16'h2A93: out_word = 8'hE6;
		16'h2A94: out_word = 8'hF1;
		16'h2A95: out_word = 8'hE3;
		16'h2A96: out_word = 8'h19;
		16'h2A97: out_word = 8'h2B;
		16'h2A98: out_word = 8'hE3;
		16'h2A99: out_word = 8'hA7;
		16'h2A9A: out_word = 8'hED;
		16'h2A9B: out_word = 8'h52;
		16'h2A9C: out_word = 8'h01;
		16'h2A9D: out_word = 8'h00;
		16'h2A9E: out_word = 8'h00;
		16'h2A9F: out_word = 8'h38;
		16'h2AA0: out_word = 8'h07;
		16'h2AA1: out_word = 8'h23;
		16'h2AA2: out_word = 8'hA7;
		16'h2AA3: out_word = 8'hFA;
		16'h2AA4: out_word = 8'h20;
		16'h2AA5: out_word = 8'h2A;
		16'h2AA6: out_word = 8'h44;
		16'h2AA7: out_word = 8'h4D;
		16'h2AA8: out_word = 8'hD1;
		16'h2AA9: out_word = 8'hFD;
		16'h2AAA: out_word = 8'hCB;
		16'h2AAB: out_word = 8'h01;
		16'h2AAC: out_word = 8'hB6;
		16'h2AAD: out_word = 8'hCD;
		16'h2AAE: out_word = 8'h30;
		16'h2AAF: out_word = 8'h25;
		16'h2AB0: out_word = 8'hC8;
		16'h2AB1: out_word = 8'hAF;
		16'h2AB2: out_word = 8'hFD;
		16'h2AB3: out_word = 8'hCB;
		16'h2AB4: out_word = 8'h01;
		16'h2AB5: out_word = 8'hB6;
		16'h2AB6: out_word = 8'hC5;
		16'h2AB7: out_word = 8'hCD;
		16'h2AB8: out_word = 8'hA9;
		16'h2AB9: out_word = 8'h33;
		16'h2ABA: out_word = 8'hC1;
		16'h2ABB: out_word = 8'h2A;
		16'h2ABC: out_word = 8'h65;
		16'h2ABD: out_word = 8'h5C;
		16'h2ABE: out_word = 8'h77;
		16'h2ABF: out_word = 8'h23;
		16'h2AC0: out_word = 8'h73;
		16'h2AC1: out_word = 8'h23;
		16'h2AC2: out_word = 8'h72;
		16'h2AC3: out_word = 8'h23;
		16'h2AC4: out_word = 8'h71;
		16'h2AC5: out_word = 8'h23;
		16'h2AC6: out_word = 8'h70;
		16'h2AC7: out_word = 8'h23;
		16'h2AC8: out_word = 8'h22;
		16'h2AC9: out_word = 8'h65;
		16'h2ACA: out_word = 8'h5C;
		16'h2ACB: out_word = 8'hC9;
		16'h2ACC: out_word = 8'hAF;
		16'h2ACD: out_word = 8'hD5;
		16'h2ACE: out_word = 8'hE5;
		16'h2ACF: out_word = 8'hF5;
		16'h2AD0: out_word = 8'hCD;
		16'h2AD1: out_word = 8'h82;
		16'h2AD2: out_word = 8'h1C;
		16'h2AD3: out_word = 8'hF1;
		16'h2AD4: out_word = 8'hCD;
		16'h2AD5: out_word = 8'h30;
		16'h2AD6: out_word = 8'h25;
		16'h2AD7: out_word = 8'h28;
		16'h2AD8: out_word = 8'h12;
		16'h2AD9: out_word = 8'hF5;
		16'h2ADA: out_word = 8'hCD;
		16'h2ADB: out_word = 8'h99;
		16'h2ADC: out_word = 8'h1E;
		16'h2ADD: out_word = 8'hD1;
		16'h2ADE: out_word = 8'h78;
		16'h2ADF: out_word = 8'hB1;
		16'h2AE0: out_word = 8'h37;
		16'h2AE1: out_word = 8'h28;
		16'h2AE2: out_word = 8'h05;
		16'h2AE3: out_word = 8'hE1;
		16'h2AE4: out_word = 8'hE5;
		16'h2AE5: out_word = 8'hA7;
		16'h2AE6: out_word = 8'hED;
		16'h2AE7: out_word = 8'h42;
		16'h2AE8: out_word = 8'h7A;
		16'h2AE9: out_word = 8'hDE;
		16'h2AEA: out_word = 8'h00;
		16'h2AEB: out_word = 8'hE1;
		16'h2AEC: out_word = 8'hD1;
		16'h2AED: out_word = 8'hC9;
		16'h2AEE: out_word = 8'hEB;
		16'h2AEF: out_word = 8'h23;
		16'h2AF0: out_word = 8'h5E;
		16'h2AF1: out_word = 8'h23;
		16'h2AF2: out_word = 8'h56;
		16'h2AF3: out_word = 8'hC9;
		16'h2AF4: out_word = 8'hCD;
		16'h2AF5: out_word = 8'h30;
		16'h2AF6: out_word = 8'h25;
		16'h2AF7: out_word = 8'hC8;
		16'h2AF8: out_word = 8'hCD;
		16'h2AF9: out_word = 8'hA9;
		16'h2AFA: out_word = 8'h30;
		16'h2AFB: out_word = 8'hDA;
		16'h2AFC: out_word = 8'h15;
		16'h2AFD: out_word = 8'h1F;
		16'h2AFE: out_word = 8'hC9;
		16'h2AFF: out_word = 8'h2A;
		16'h2B00: out_word = 8'h4D;
		16'h2B01: out_word = 8'h5C;
		16'h2B02: out_word = 8'hFD;
		16'h2B03: out_word = 8'hCB;
		16'h2B04: out_word = 8'h37;
		16'h2B05: out_word = 8'h4E;
		16'h2B06: out_word = 8'h28;
		16'h2B07: out_word = 8'h5E;
		16'h2B08: out_word = 8'h01;
		16'h2B09: out_word = 8'h05;
		16'h2B0A: out_word = 8'h00;
		16'h2B0B: out_word = 8'h03;
		16'h2B0C: out_word = 8'h23;
		16'h2B0D: out_word = 8'h7E;
		16'h2B0E: out_word = 8'hFE;
		16'h2B0F: out_word = 8'h20;
		16'h2B10: out_word = 8'h28;
		16'h2B11: out_word = 8'hFA;
		16'h2B12: out_word = 8'h30;
		16'h2B13: out_word = 8'h0B;
		16'h2B14: out_word = 8'hFE;
		16'h2B15: out_word = 8'h10;
		16'h2B16: out_word = 8'h38;
		16'h2B17: out_word = 8'h11;
		16'h2B18: out_word = 8'hFE;
		16'h2B19: out_word = 8'h16;
		16'h2B1A: out_word = 8'h30;
		16'h2B1B: out_word = 8'h0D;
		16'h2B1C: out_word = 8'h23;
		16'h2B1D: out_word = 8'h18;
		16'h2B1E: out_word = 8'hED;
		16'h2B1F: out_word = 8'hCD;
		16'h2B20: out_word = 8'h88;
		16'h2B21: out_word = 8'h2C;
		16'h2B22: out_word = 8'h38;
		16'h2B23: out_word = 8'hE7;
		16'h2B24: out_word = 8'hFE;
		16'h2B25: out_word = 8'h24;
		16'h2B26: out_word = 8'hCA;
		16'h2B27: out_word = 8'hC0;
		16'h2B28: out_word = 8'h2B;
		16'h2B29: out_word = 8'h79;
		16'h2B2A: out_word = 8'h2A;
		16'h2B2B: out_word = 8'h59;
		16'h2B2C: out_word = 8'h5C;
		16'h2B2D: out_word = 8'h2B;
		16'h2B2E: out_word = 8'hCD;
		16'h2B2F: out_word = 8'h55;
		16'h2B30: out_word = 8'h16;
		16'h2B31: out_word = 8'h23;
		16'h2B32: out_word = 8'h23;
		16'h2B33: out_word = 8'hEB;
		16'h2B34: out_word = 8'hD5;
		16'h2B35: out_word = 8'h2A;
		16'h2B36: out_word = 8'h4D;
		16'h2B37: out_word = 8'h5C;
		16'h2B38: out_word = 8'h1B;
		16'h2B39: out_word = 8'hD6;
		16'h2B3A: out_word = 8'h06;
		16'h2B3B: out_word = 8'h47;
		16'h2B3C: out_word = 8'h28;
		16'h2B3D: out_word = 8'h11;
		16'h2B3E: out_word = 8'h23;
		16'h2B3F: out_word = 8'h7E;
		16'h2B40: out_word = 8'hFE;
		16'h2B41: out_word = 8'h21;
		16'h2B42: out_word = 8'h38;
		16'h2B43: out_word = 8'hFA;
		16'h2B44: out_word = 8'hF6;
		16'h2B45: out_word = 8'h20;
		16'h2B46: out_word = 8'h13;
		16'h2B47: out_word = 8'h12;
		16'h2B48: out_word = 8'h10;
		16'h2B49: out_word = 8'hF4;
		16'h2B4A: out_word = 8'hF6;
		16'h2B4B: out_word = 8'h80;
		16'h2B4C: out_word = 8'h12;
		16'h2B4D: out_word = 8'h3E;
		16'h2B4E: out_word = 8'hC0;
		16'h2B4F: out_word = 8'h2A;
		16'h2B50: out_word = 8'h4D;
		16'h2B51: out_word = 8'h5C;
		16'h2B52: out_word = 8'hAE;
		16'h2B53: out_word = 8'hF6;
		16'h2B54: out_word = 8'h20;
		16'h2B55: out_word = 8'hE1;
		16'h2B56: out_word = 8'hCD;
		16'h2B57: out_word = 8'hEA;
		16'h2B58: out_word = 8'h2B;
		16'h2B59: out_word = 8'hE5;
		16'h2B5A: out_word = 8'hEF;
		16'h2B5B: out_word = 8'h02;
		16'h2B5C: out_word = 8'h38;
		16'h2B5D: out_word = 8'hE1;
		16'h2B5E: out_word = 8'h01;
		16'h2B5F: out_word = 8'h05;
		16'h2B60: out_word = 8'h00;
		16'h2B61: out_word = 8'hA7;
		16'h2B62: out_word = 8'hED;
		16'h2B63: out_word = 8'h42;
		16'h2B64: out_word = 8'h18;
		16'h2B65: out_word = 8'h40;
		16'h2B66: out_word = 8'hFD;
		16'h2B67: out_word = 8'hCB;
		16'h2B68: out_word = 8'h01;
		16'h2B69: out_word = 8'h76;
		16'h2B6A: out_word = 8'h28;
		16'h2B6B: out_word = 8'h06;
		16'h2B6C: out_word = 8'h11;
		16'h2B6D: out_word = 8'h06;
		16'h2B6E: out_word = 8'h00;
		16'h2B6F: out_word = 8'h19;
		16'h2B70: out_word = 8'h18;
		16'h2B71: out_word = 8'hE7;
		16'h2B72: out_word = 8'h2A;
		16'h2B73: out_word = 8'h4D;
		16'h2B74: out_word = 8'h5C;
		16'h2B75: out_word = 8'hED;
		16'h2B76: out_word = 8'h4B;
		16'h2B77: out_word = 8'h72;
		16'h2B78: out_word = 8'h5C;
		16'h2B79: out_word = 8'hFD;
		16'h2B7A: out_word = 8'hCB;
		16'h2B7B: out_word = 8'h37;
		16'h2B7C: out_word = 8'h46;
		16'h2B7D: out_word = 8'h20;
		16'h2B7E: out_word = 8'h30;
		16'h2B7F: out_word = 8'h78;
		16'h2B80: out_word = 8'hB1;
		16'h2B81: out_word = 8'hC8;
		16'h2B82: out_word = 8'hE5;
		16'h2B83: out_word = 8'hF7;
		16'h2B84: out_word = 8'hD5;
		16'h2B85: out_word = 8'hC5;
		16'h2B86: out_word = 8'h54;
		16'h2B87: out_word = 8'h5D;
		16'h2B88: out_word = 8'h23;
		16'h2B89: out_word = 8'h36;
		16'h2B8A: out_word = 8'h20;
		16'h2B8B: out_word = 8'hED;
		16'h2B8C: out_word = 8'hB8;
		16'h2B8D: out_word = 8'hE5;
		16'h2B8E: out_word = 8'hCD;
		16'h2B8F: out_word = 8'hF1;
		16'h2B90: out_word = 8'h2B;
		16'h2B91: out_word = 8'hE1;
		16'h2B92: out_word = 8'hE3;
		16'h2B93: out_word = 8'hA7;
		16'h2B94: out_word = 8'hED;
		16'h2B95: out_word = 8'h42;
		16'h2B96: out_word = 8'h09;
		16'h2B97: out_word = 8'h30;
		16'h2B98: out_word = 8'h02;
		16'h2B99: out_word = 8'h44;
		16'h2B9A: out_word = 8'h4D;
		16'h2B9B: out_word = 8'hE3;
		16'h2B9C: out_word = 8'hEB;
		16'h2B9D: out_word = 8'h78;
		16'h2B9E: out_word = 8'hB1;
		16'h2B9F: out_word = 8'h28;
		16'h2BA0: out_word = 8'h02;
		16'h2BA1: out_word = 8'hED;
		16'h2BA2: out_word = 8'hB0;
		16'h2BA3: out_word = 8'hC1;
		16'h2BA4: out_word = 8'hD1;
		16'h2BA5: out_word = 8'hE1;
		16'h2BA6: out_word = 8'hEB;
		16'h2BA7: out_word = 8'h78;
		16'h2BA8: out_word = 8'hB1;
		16'h2BA9: out_word = 8'hC8;
		16'h2BAA: out_word = 8'hD5;
		16'h2BAB: out_word = 8'hED;
		16'h2BAC: out_word = 8'hB0;
		16'h2BAD: out_word = 8'hE1;
		16'h2BAE: out_word = 8'hC9;
		16'h2BAF: out_word = 8'h2B;
		16'h2BB0: out_word = 8'h2B;
		16'h2BB1: out_word = 8'h2B;
		16'h2BB2: out_word = 8'h7E;
		16'h2BB3: out_word = 8'hE5;
		16'h2BB4: out_word = 8'hC5;
		16'h2BB5: out_word = 8'hCD;
		16'h2BB6: out_word = 8'hC6;
		16'h2BB7: out_word = 8'h2B;
		16'h2BB8: out_word = 8'hC1;
		16'h2BB9: out_word = 8'hE1;
		16'h2BBA: out_word = 8'h03;
		16'h2BBB: out_word = 8'h03;
		16'h2BBC: out_word = 8'h03;
		16'h2BBD: out_word = 8'hC3;
		16'h2BBE: out_word = 8'hE8;
		16'h2BBF: out_word = 8'h19;
		16'h2BC0: out_word = 8'h3E;
		16'h2BC1: out_word = 8'hDF;
		16'h2BC2: out_word = 8'h2A;
		16'h2BC3: out_word = 8'h4D;
		16'h2BC4: out_word = 8'h5C;
		16'h2BC5: out_word = 8'hA6;
		16'h2BC6: out_word = 8'hF5;
		16'h2BC7: out_word = 8'hCD;
		16'h2BC8: out_word = 8'hF1;
		16'h2BC9: out_word = 8'h2B;
		16'h2BCA: out_word = 8'hEB;
		16'h2BCB: out_word = 8'h09;
		16'h2BCC: out_word = 8'hC5;
		16'h2BCD: out_word = 8'h2B;
		16'h2BCE: out_word = 8'h22;
		16'h2BCF: out_word = 8'h4D;
		16'h2BD0: out_word = 8'h5C;
		16'h2BD1: out_word = 8'h03;
		16'h2BD2: out_word = 8'h03;
		16'h2BD3: out_word = 8'h03;
		16'h2BD4: out_word = 8'h2A;
		16'h2BD5: out_word = 8'h59;
		16'h2BD6: out_word = 8'h5C;
		16'h2BD7: out_word = 8'h2B;
		16'h2BD8: out_word = 8'hCD;
		16'h2BD9: out_word = 8'h55;
		16'h2BDA: out_word = 8'h16;
		16'h2BDB: out_word = 8'h2A;
		16'h2BDC: out_word = 8'h4D;
		16'h2BDD: out_word = 8'h5C;
		16'h2BDE: out_word = 8'hC1;
		16'h2BDF: out_word = 8'hC5;
		16'h2BE0: out_word = 8'h03;
		16'h2BE1: out_word = 8'hED;
		16'h2BE2: out_word = 8'hB8;
		16'h2BE3: out_word = 8'hEB;
		16'h2BE4: out_word = 8'h23;
		16'h2BE5: out_word = 8'hC1;
		16'h2BE6: out_word = 8'h70;
		16'h2BE7: out_word = 8'h2B;
		16'h2BE8: out_word = 8'h71;
		16'h2BE9: out_word = 8'hF1;
		16'h2BEA: out_word = 8'h2B;
		16'h2BEB: out_word = 8'h77;
		16'h2BEC: out_word = 8'h2A;
		16'h2BED: out_word = 8'h59;
		16'h2BEE: out_word = 8'h5C;
		16'h2BEF: out_word = 8'h2B;
		16'h2BF0: out_word = 8'hC9;
		16'h2BF1: out_word = 8'h2A;
		16'h2BF2: out_word = 8'h65;
		16'h2BF3: out_word = 8'h5C;
		16'h2BF4: out_word = 8'h2B;
		16'h2BF5: out_word = 8'h46;
		16'h2BF6: out_word = 8'h2B;
		16'h2BF7: out_word = 8'h4E;
		16'h2BF8: out_word = 8'h2B;
		16'h2BF9: out_word = 8'h56;
		16'h2BFA: out_word = 8'h2B;
		16'h2BFB: out_word = 8'h5E;
		16'h2BFC: out_word = 8'h2B;
		16'h2BFD: out_word = 8'h7E;
		16'h2BFE: out_word = 8'h22;
		16'h2BFF: out_word = 8'h65;
		16'h2C00: out_word = 8'h5C;
		16'h2C01: out_word = 8'hC9;
		16'h2C02: out_word = 8'hCD;
		16'h2C03: out_word = 8'hB2;
		16'h2C04: out_word = 8'h28;
		16'h2C05: out_word = 8'hC2;
		16'h2C06: out_word = 8'h8A;
		16'h2C07: out_word = 8'h1C;
		16'h2C08: out_word = 8'hCD;
		16'h2C09: out_word = 8'h30;
		16'h2C0A: out_word = 8'h25;
		16'h2C0B: out_word = 8'h20;
		16'h2C0C: out_word = 8'h08;
		16'h2C0D: out_word = 8'hCB;
		16'h2C0E: out_word = 8'hB1;
		16'h2C0F: out_word = 8'hCD;
		16'h2C10: out_word = 8'h96;
		16'h2C11: out_word = 8'h29;
		16'h2C12: out_word = 8'hCD;
		16'h2C13: out_word = 8'hEE;
		16'h2C14: out_word = 8'h1B;
		16'h2C15: out_word = 8'h38;
		16'h2C16: out_word = 8'h08;
		16'h2C17: out_word = 8'hC5;
		16'h2C18: out_word = 8'hCD;
		16'h2C19: out_word = 8'hB8;
		16'h2C1A: out_word = 8'h19;
		16'h2C1B: out_word = 8'hCD;
		16'h2C1C: out_word = 8'hE8;
		16'h2C1D: out_word = 8'h19;
		16'h2C1E: out_word = 8'hC1;
		16'h2C1F: out_word = 8'hCB;
		16'h2C20: out_word = 8'hF9;
		16'h2C21: out_word = 8'h06;
		16'h2C22: out_word = 8'h00;
		16'h2C23: out_word = 8'hC5;
		16'h2C24: out_word = 8'h21;
		16'h2C25: out_word = 8'h01;
		16'h2C26: out_word = 8'h00;
		16'h2C27: out_word = 8'hCB;
		16'h2C28: out_word = 8'h71;
		16'h2C29: out_word = 8'h20;
		16'h2C2A: out_word = 8'h02;
		16'h2C2B: out_word = 8'h2E;
		16'h2C2C: out_word = 8'h05;
		16'h2C2D: out_word = 8'hEB;
		16'h2C2E: out_word = 8'hE7;
		16'h2C2F: out_word = 8'h26;
		16'h2C30: out_word = 8'hFF;
		16'h2C31: out_word = 8'hCD;
		16'h2C32: out_word = 8'hCC;
		16'h2C33: out_word = 8'h2A;
		16'h2C34: out_word = 8'hDA;
		16'h2C35: out_word = 8'h20;
		16'h2C36: out_word = 8'h2A;
		16'h2C37: out_word = 8'hE1;
		16'h2C38: out_word = 8'hC5;
		16'h2C39: out_word = 8'h24;
		16'h2C3A: out_word = 8'hE5;
		16'h2C3B: out_word = 8'h60;
		16'h2C3C: out_word = 8'h69;
		16'h2C3D: out_word = 8'hCD;
		16'h2C3E: out_word = 8'hF4;
		16'h2C3F: out_word = 8'h2A;
		16'h2C40: out_word = 8'hEB;
		16'h2C41: out_word = 8'hDF;
		16'h2C42: out_word = 8'hFE;
		16'h2C43: out_word = 8'h2C;
		16'h2C44: out_word = 8'h28;
		16'h2C45: out_word = 8'hE8;
		16'h2C46: out_word = 8'hFE;
		16'h2C47: out_word = 8'h29;
		16'h2C48: out_word = 8'h20;
		16'h2C49: out_word = 8'hBB;
		16'h2C4A: out_word = 8'hE7;
		16'h2C4B: out_word = 8'hC1;
		16'h2C4C: out_word = 8'h79;
		16'h2C4D: out_word = 8'h68;
		16'h2C4E: out_word = 8'h26;
		16'h2C4F: out_word = 8'h00;
		16'h2C50: out_word = 8'h23;
		16'h2C51: out_word = 8'h23;
		16'h2C52: out_word = 8'h29;
		16'h2C53: out_word = 8'h19;
		16'h2C54: out_word = 8'hDA;
		16'h2C55: out_word = 8'h15;
		16'h2C56: out_word = 8'h1F;
		16'h2C57: out_word = 8'hD5;
		16'h2C58: out_word = 8'hC5;
		16'h2C59: out_word = 8'hE5;
		16'h2C5A: out_word = 8'h44;
		16'h2C5B: out_word = 8'h4D;
		16'h2C5C: out_word = 8'h2A;
		16'h2C5D: out_word = 8'h59;
		16'h2C5E: out_word = 8'h5C;
		16'h2C5F: out_word = 8'h2B;
		16'h2C60: out_word = 8'hCD;
		16'h2C61: out_word = 8'h55;
		16'h2C62: out_word = 8'h16;
		16'h2C63: out_word = 8'h23;
		16'h2C64: out_word = 8'h77;
		16'h2C65: out_word = 8'hC1;
		16'h2C66: out_word = 8'h0B;
		16'h2C67: out_word = 8'h0B;
		16'h2C68: out_word = 8'h0B;
		16'h2C69: out_word = 8'h23;
		16'h2C6A: out_word = 8'h71;
		16'h2C6B: out_word = 8'h23;
		16'h2C6C: out_word = 8'h70;
		16'h2C6D: out_word = 8'hC1;
		16'h2C6E: out_word = 8'h78;
		16'h2C6F: out_word = 8'h23;
		16'h2C70: out_word = 8'h77;
		16'h2C71: out_word = 8'h62;
		16'h2C72: out_word = 8'h6B;
		16'h2C73: out_word = 8'h1B;
		16'h2C74: out_word = 8'h36;
		16'h2C75: out_word = 8'h00;
		16'h2C76: out_word = 8'hCB;
		16'h2C77: out_word = 8'h71;
		16'h2C78: out_word = 8'h28;
		16'h2C79: out_word = 8'h02;
		16'h2C7A: out_word = 8'h36;
		16'h2C7B: out_word = 8'h20;
		16'h2C7C: out_word = 8'hC1;
		16'h2C7D: out_word = 8'hED;
		16'h2C7E: out_word = 8'hB8;
		16'h2C7F: out_word = 8'hC1;
		16'h2C80: out_word = 8'h70;
		16'h2C81: out_word = 8'h2B;
		16'h2C82: out_word = 8'h71;
		16'h2C83: out_word = 8'h2B;
		16'h2C84: out_word = 8'h3D;
		16'h2C85: out_word = 8'h20;
		16'h2C86: out_word = 8'hF8;
		16'h2C87: out_word = 8'hC9;
		16'h2C88: out_word = 8'hCD;
		16'h2C89: out_word = 8'h1B;
		16'h2C8A: out_word = 8'h2D;
		16'h2C8B: out_word = 8'h3F;
		16'h2C8C: out_word = 8'hD8;
		16'h2C8D: out_word = 8'hFE;
		16'h2C8E: out_word = 8'h41;
		16'h2C8F: out_word = 8'h3F;
		16'h2C90: out_word = 8'hD0;
		16'h2C91: out_word = 8'hFE;
		16'h2C92: out_word = 8'h5B;
		16'h2C93: out_word = 8'hD8;
		16'h2C94: out_word = 8'hFE;
		16'h2C95: out_word = 8'h61;
		16'h2C96: out_word = 8'h3F;
		16'h2C97: out_word = 8'hD0;
		16'h2C98: out_word = 8'hFE;
		16'h2C99: out_word = 8'h7B;
		16'h2C9A: out_word = 8'hC9;
		16'h2C9B: out_word = 8'hFE;
		16'h2C9C: out_word = 8'hC4;
		16'h2C9D: out_word = 8'h20;
		16'h2C9E: out_word = 8'h19;
		16'h2C9F: out_word = 8'h11;
		16'h2CA0: out_word = 8'h00;
		16'h2CA1: out_word = 8'h00;
		16'h2CA2: out_word = 8'hE7;
		16'h2CA3: out_word = 8'hD6;
		16'h2CA4: out_word = 8'h31;
		16'h2CA5: out_word = 8'hCE;
		16'h2CA6: out_word = 8'h00;
		16'h2CA7: out_word = 8'h20;
		16'h2CA8: out_word = 8'h0A;
		16'h2CA9: out_word = 8'hEB;
		16'h2CAA: out_word = 8'h3F;
		16'h2CAB: out_word = 8'hED;
		16'h2CAC: out_word = 8'h6A;
		16'h2CAD: out_word = 8'hDA;
		16'h2CAE: out_word = 8'hAD;
		16'h2CAF: out_word = 8'h31;
		16'h2CB0: out_word = 8'hEB;
		16'h2CB1: out_word = 8'h18;
		16'h2CB2: out_word = 8'hEF;
		16'h2CB3: out_word = 8'h42;
		16'h2CB4: out_word = 8'h4B;
		16'h2CB5: out_word = 8'hC3;
		16'h2CB6: out_word = 8'h2B;
		16'h2CB7: out_word = 8'h2D;
		16'h2CB8: out_word = 8'hFE;
		16'h2CB9: out_word = 8'h2E;
		16'h2CBA: out_word = 8'h28;
		16'h2CBB: out_word = 8'h0F;
		16'h2CBC: out_word = 8'hCD;
		16'h2CBD: out_word = 8'h3B;
		16'h2CBE: out_word = 8'h2D;
		16'h2CBF: out_word = 8'hFE;
		16'h2CC0: out_word = 8'h2E;
		16'h2CC1: out_word = 8'h20;
		16'h2CC2: out_word = 8'h28;
		16'h2CC3: out_word = 8'hE7;
		16'h2CC4: out_word = 8'hCD;
		16'h2CC5: out_word = 8'h1B;
		16'h2CC6: out_word = 8'h2D;
		16'h2CC7: out_word = 8'h38;
		16'h2CC8: out_word = 8'h22;
		16'h2CC9: out_word = 8'h18;
		16'h2CCA: out_word = 8'h0A;
		16'h2CCB: out_word = 8'hE7;
		16'h2CCC: out_word = 8'hCD;
		16'h2CCD: out_word = 8'h1B;
		16'h2CCE: out_word = 8'h2D;
		16'h2CCF: out_word = 8'hDA;
		16'h2CD0: out_word = 8'h8A;
		16'h2CD1: out_word = 8'h1C;
		16'h2CD2: out_word = 8'hEF;
		16'h2CD3: out_word = 8'hA0;
		16'h2CD4: out_word = 8'h38;
		16'h2CD5: out_word = 8'hEF;
		16'h2CD6: out_word = 8'hA1;
		16'h2CD7: out_word = 8'hC0;
		16'h2CD8: out_word = 8'h02;
		16'h2CD9: out_word = 8'h38;
		16'h2CDA: out_word = 8'hDF;
		16'h2CDB: out_word = 8'hCD;
		16'h2CDC: out_word = 8'h22;
		16'h2CDD: out_word = 8'h2D;
		16'h2CDE: out_word = 8'h38;
		16'h2CDF: out_word = 8'h0B;
		16'h2CE0: out_word = 8'hEF;
		16'h2CE1: out_word = 8'hE0;
		16'h2CE2: out_word = 8'hA4;
		16'h2CE3: out_word = 8'h05;
		16'h2CE4: out_word = 8'hC0;
		16'h2CE5: out_word = 8'h04;
		16'h2CE6: out_word = 8'h0F;
		16'h2CE7: out_word = 8'h38;
		16'h2CE8: out_word = 8'hE7;
		16'h2CE9: out_word = 8'h18;
		16'h2CEA: out_word = 8'hEF;
		16'h2CEB: out_word = 8'hFE;
		16'h2CEC: out_word = 8'h45;
		16'h2CED: out_word = 8'h28;
		16'h2CEE: out_word = 8'h03;
		16'h2CEF: out_word = 8'hFE;
		16'h2CF0: out_word = 8'h65;
		16'h2CF1: out_word = 8'hC0;
		16'h2CF2: out_word = 8'h06;
		16'h2CF3: out_word = 8'hFF;
		16'h2CF4: out_word = 8'hE7;
		16'h2CF5: out_word = 8'hFE;
		16'h2CF6: out_word = 8'h2B;
		16'h2CF7: out_word = 8'h28;
		16'h2CF8: out_word = 8'h05;
		16'h2CF9: out_word = 8'hFE;
		16'h2CFA: out_word = 8'h2D;
		16'h2CFB: out_word = 8'h20;
		16'h2CFC: out_word = 8'h02;
		16'h2CFD: out_word = 8'h04;
		16'h2CFE: out_word = 8'hE7;
		16'h2CFF: out_word = 8'hCD;
		16'h2D00: out_word = 8'h1B;
		16'h2D01: out_word = 8'h2D;
		16'h2D02: out_word = 8'h38;
		16'h2D03: out_word = 8'hCB;
		16'h2D04: out_word = 8'hC5;
		16'h2D05: out_word = 8'hCD;
		16'h2D06: out_word = 8'h3B;
		16'h2D07: out_word = 8'h2D;
		16'h2D08: out_word = 8'hCD;
		16'h2D09: out_word = 8'hD5;
		16'h2D0A: out_word = 8'h2D;
		16'h2D0B: out_word = 8'hC1;
		16'h2D0C: out_word = 8'hDA;
		16'h2D0D: out_word = 8'hAD;
		16'h2D0E: out_word = 8'h31;
		16'h2D0F: out_word = 8'hA7;
		16'h2D10: out_word = 8'hFA;
		16'h2D11: out_word = 8'hAD;
		16'h2D12: out_word = 8'h31;
		16'h2D13: out_word = 8'h04;
		16'h2D14: out_word = 8'h28;
		16'h2D15: out_word = 8'h02;
		16'h2D16: out_word = 8'hED;
		16'h2D17: out_word = 8'h44;
		16'h2D18: out_word = 8'hC3;
		16'h2D19: out_word = 8'h4F;
		16'h2D1A: out_word = 8'h2D;
		16'h2D1B: out_word = 8'hFE;
		16'h2D1C: out_word = 8'h30;
		16'h2D1D: out_word = 8'hD8;
		16'h2D1E: out_word = 8'hFE;
		16'h2D1F: out_word = 8'h3A;
		16'h2D20: out_word = 8'h3F;
		16'h2D21: out_word = 8'hC9;
		16'h2D22: out_word = 8'hCD;
		16'h2D23: out_word = 8'h1B;
		16'h2D24: out_word = 8'h2D;
		16'h2D25: out_word = 8'hD8;
		16'h2D26: out_word = 8'hD6;
		16'h2D27: out_word = 8'h30;
		16'h2D28: out_word = 8'h4F;
		16'h2D29: out_word = 8'h06;
		16'h2D2A: out_word = 8'h00;
		16'h2D2B: out_word = 8'hFD;
		16'h2D2C: out_word = 8'h21;
		16'h2D2D: out_word = 8'h3A;
		16'h2D2E: out_word = 8'h5C;
		16'h2D2F: out_word = 8'hAF;
		16'h2D30: out_word = 8'h5F;
		16'h2D31: out_word = 8'h51;
		16'h2D32: out_word = 8'h48;
		16'h2D33: out_word = 8'h47;
		16'h2D34: out_word = 8'hCD;
		16'h2D35: out_word = 8'hB6;
		16'h2D36: out_word = 8'h2A;
		16'h2D37: out_word = 8'hEF;
		16'h2D38: out_word = 8'h38;
		16'h2D39: out_word = 8'hA7;
		16'h2D3A: out_word = 8'hC9;
		16'h2D3B: out_word = 8'hF5;
		16'h2D3C: out_word = 8'hEF;
		16'h2D3D: out_word = 8'hA0;
		16'h2D3E: out_word = 8'h38;
		16'h2D3F: out_word = 8'hF1;
		16'h2D40: out_word = 8'hCD;
		16'h2D41: out_word = 8'h22;
		16'h2D42: out_word = 8'h2D;
		16'h2D43: out_word = 8'hD8;
		16'h2D44: out_word = 8'hEF;
		16'h2D45: out_word = 8'h01;
		16'h2D46: out_word = 8'hA4;
		16'h2D47: out_word = 8'h04;
		16'h2D48: out_word = 8'h0F;
		16'h2D49: out_word = 8'h38;
		16'h2D4A: out_word = 8'hCD;
		16'h2D4B: out_word = 8'h74;
		16'h2D4C: out_word = 8'h00;
		16'h2D4D: out_word = 8'h18;
		16'h2D4E: out_word = 8'hF1;
		16'h2D4F: out_word = 8'h07;
		16'h2D50: out_word = 8'h0F;
		16'h2D51: out_word = 8'h30;
		16'h2D52: out_word = 8'h02;
		16'h2D53: out_word = 8'h2F;
		16'h2D54: out_word = 8'h3C;
		16'h2D55: out_word = 8'hF5;
		16'h2D56: out_word = 8'h21;
		16'h2D57: out_word = 8'h92;
		16'h2D58: out_word = 8'h5C;
		16'h2D59: out_word = 8'hCD;
		16'h2D5A: out_word = 8'h0B;
		16'h2D5B: out_word = 8'h35;
		16'h2D5C: out_word = 8'hEF;
		16'h2D5D: out_word = 8'hA4;
		16'h2D5E: out_word = 8'h38;
		16'h2D5F: out_word = 8'hF1;
		16'h2D60: out_word = 8'hCB;
		16'h2D61: out_word = 8'h3F;
		16'h2D62: out_word = 8'h30;
		16'h2D63: out_word = 8'h0D;
		16'h2D64: out_word = 8'hF5;
		16'h2D65: out_word = 8'hEF;
		16'h2D66: out_word = 8'hC1;
		16'h2D67: out_word = 8'hE0;
		16'h2D68: out_word = 8'h00;
		16'h2D69: out_word = 8'h04;
		16'h2D6A: out_word = 8'h04;
		16'h2D6B: out_word = 8'h33;
		16'h2D6C: out_word = 8'h02;
		16'h2D6D: out_word = 8'h05;
		16'h2D6E: out_word = 8'hE1;
		16'h2D6F: out_word = 8'h38;
		16'h2D70: out_word = 8'hF1;
		16'h2D71: out_word = 8'h28;
		16'h2D72: out_word = 8'h08;
		16'h2D73: out_word = 8'hF5;
		16'h2D74: out_word = 8'hEF;
		16'h2D75: out_word = 8'h31;
		16'h2D76: out_word = 8'h04;
		16'h2D77: out_word = 8'h38;
		16'h2D78: out_word = 8'hF1;
		16'h2D79: out_word = 8'h18;
		16'h2D7A: out_word = 8'hE5;
		16'h2D7B: out_word = 8'hEF;
		16'h2D7C: out_word = 8'h02;
		16'h2D7D: out_word = 8'h38;
		16'h2D7E: out_word = 8'hC9;
		16'h2D7F: out_word = 8'h23;
		16'h2D80: out_word = 8'h4E;
		16'h2D81: out_word = 8'h23;
		16'h2D82: out_word = 8'h7E;
		16'h2D83: out_word = 8'hA9;
		16'h2D84: out_word = 8'h91;
		16'h2D85: out_word = 8'h5F;
		16'h2D86: out_word = 8'h23;
		16'h2D87: out_word = 8'h7E;
		16'h2D88: out_word = 8'h89;
		16'h2D89: out_word = 8'hA9;
		16'h2D8A: out_word = 8'h57;
		16'h2D8B: out_word = 8'hC9;
		16'h2D8C: out_word = 8'h0E;
		16'h2D8D: out_word = 8'h00;
		16'h2D8E: out_word = 8'hE5;
		16'h2D8F: out_word = 8'h36;
		16'h2D90: out_word = 8'h00;
		16'h2D91: out_word = 8'h23;
		16'h2D92: out_word = 8'h71;
		16'h2D93: out_word = 8'h23;
		16'h2D94: out_word = 8'h7B;
		16'h2D95: out_word = 8'hA9;
		16'h2D96: out_word = 8'h91;
		16'h2D97: out_word = 8'h77;
		16'h2D98: out_word = 8'h23;
		16'h2D99: out_word = 8'h7A;
		16'h2D9A: out_word = 8'h89;
		16'h2D9B: out_word = 8'hA9;
		16'h2D9C: out_word = 8'h77;
		16'h2D9D: out_word = 8'h23;
		16'h2D9E: out_word = 8'h36;
		16'h2D9F: out_word = 8'h00;
		16'h2DA0: out_word = 8'hE1;
		16'h2DA1: out_word = 8'hC9;
		16'h2DA2: out_word = 8'hEF;
		16'h2DA3: out_word = 8'h38;
		16'h2DA4: out_word = 8'h7E;
		16'h2DA5: out_word = 8'hA7;
		16'h2DA6: out_word = 8'h28;
		16'h2DA7: out_word = 8'h05;
		16'h2DA8: out_word = 8'hEF;
		16'h2DA9: out_word = 8'hA2;
		16'h2DAA: out_word = 8'h0F;
		16'h2DAB: out_word = 8'h27;
		16'h2DAC: out_word = 8'h38;
		16'h2DAD: out_word = 8'hEF;
		16'h2DAE: out_word = 8'h02;
		16'h2DAF: out_word = 8'h38;
		16'h2DB0: out_word = 8'hE5;
		16'h2DB1: out_word = 8'hD5;
		16'h2DB2: out_word = 8'hEB;
		16'h2DB3: out_word = 8'h46;
		16'h2DB4: out_word = 8'hCD;
		16'h2DB5: out_word = 8'h7F;
		16'h2DB6: out_word = 8'h2D;
		16'h2DB7: out_word = 8'hAF;
		16'h2DB8: out_word = 8'h90;
		16'h2DB9: out_word = 8'hCB;
		16'h2DBA: out_word = 8'h79;
		16'h2DBB: out_word = 8'h42;
		16'h2DBC: out_word = 8'h4B;
		16'h2DBD: out_word = 8'h7B;
		16'h2DBE: out_word = 8'hD1;
		16'h2DBF: out_word = 8'hE1;
		16'h2DC0: out_word = 8'hC9;
		16'h2DC1: out_word = 8'h57;
		16'h2DC2: out_word = 8'h17;
		16'h2DC3: out_word = 8'h9F;
		16'h2DC4: out_word = 8'h5F;
		16'h2DC5: out_word = 8'h4F;
		16'h2DC6: out_word = 8'hAF;
		16'h2DC7: out_word = 8'h47;
		16'h2DC8: out_word = 8'hCD;
		16'h2DC9: out_word = 8'hB6;
		16'h2DCA: out_word = 8'h2A;
		16'h2DCB: out_word = 8'hEF;
		16'h2DCC: out_word = 8'h34;
		16'h2DCD: out_word = 8'hEF;
		16'h2DCE: out_word = 8'h1A;
		16'h2DCF: out_word = 8'h20;
		16'h2DD0: out_word = 8'h9A;
		16'h2DD1: out_word = 8'h85;
		16'h2DD2: out_word = 8'h04;
		16'h2DD3: out_word = 8'h27;
		16'h2DD4: out_word = 8'h38;
		16'h2DD5: out_word = 8'hCD;
		16'h2DD6: out_word = 8'hA2;
		16'h2DD7: out_word = 8'h2D;
		16'h2DD8: out_word = 8'hD8;
		16'h2DD9: out_word = 8'hF5;
		16'h2DDA: out_word = 8'h05;
		16'h2DDB: out_word = 8'h04;
		16'h2DDC: out_word = 8'h28;
		16'h2DDD: out_word = 8'h03;
		16'h2DDE: out_word = 8'hF1;
		16'h2DDF: out_word = 8'h37;
		16'h2DE0: out_word = 8'hC9;
		16'h2DE1: out_word = 8'hF1;
		16'h2DE2: out_word = 8'hC9;
		16'h2DE3: out_word = 8'hEF;
		16'h2DE4: out_word = 8'h31;
		16'h2DE5: out_word = 8'h36;
		16'h2DE6: out_word = 8'h00;
		16'h2DE7: out_word = 8'h0B;
		16'h2DE8: out_word = 8'h31;
		16'h2DE9: out_word = 8'h37;
		16'h2DEA: out_word = 8'h00;
		16'h2DEB: out_word = 8'h0D;
		16'h2DEC: out_word = 8'h02;
		16'h2DED: out_word = 8'h38;
		16'h2DEE: out_word = 8'h3E;
		16'h2DEF: out_word = 8'h30;
		16'h2DF0: out_word = 8'hD7;
		16'h2DF1: out_word = 8'hC9;
		16'h2DF2: out_word = 8'h2A;
		16'h2DF3: out_word = 8'h38;
		16'h2DF4: out_word = 8'h3E;
		16'h2DF5: out_word = 8'h2D;
		16'h2DF6: out_word = 8'hD7;
		16'h2DF7: out_word = 8'hEF;
		16'h2DF8: out_word = 8'hA0;
		16'h2DF9: out_word = 8'hC3;
		16'h2DFA: out_word = 8'hC4;
		16'h2DFB: out_word = 8'hC5;
		16'h2DFC: out_word = 8'h02;
		16'h2DFD: out_word = 8'h38;
		16'h2DFE: out_word = 8'hD9;
		16'h2DFF: out_word = 8'hE5;
		16'h2E00: out_word = 8'hD9;
		16'h2E01: out_word = 8'hEF;
		16'h2E02: out_word = 8'h31;
		16'h2E03: out_word = 8'h27;
		16'h2E04: out_word = 8'hC2;
		16'h2E05: out_word = 8'h03;
		16'h2E06: out_word = 8'hE2;
		16'h2E07: out_word = 8'h01;
		16'h2E08: out_word = 8'hC2;
		16'h2E09: out_word = 8'h02;
		16'h2E0A: out_word = 8'h38;
		16'h2E0B: out_word = 8'h7E;
		16'h2E0C: out_word = 8'hA7;
		16'h2E0D: out_word = 8'h20;
		16'h2E0E: out_word = 8'h47;
		16'h2E0F: out_word = 8'hCD;
		16'h2E10: out_word = 8'h7F;
		16'h2E11: out_word = 8'h2D;
		16'h2E12: out_word = 8'h06;
		16'h2E13: out_word = 8'h10;
		16'h2E14: out_word = 8'h7A;
		16'h2E15: out_word = 8'hA7;
		16'h2E16: out_word = 8'h20;
		16'h2E17: out_word = 8'h06;
		16'h2E18: out_word = 8'hB3;
		16'h2E19: out_word = 8'h28;
		16'h2E1A: out_word = 8'h09;
		16'h2E1B: out_word = 8'h53;
		16'h2E1C: out_word = 8'h06;
		16'h2E1D: out_word = 8'h08;
		16'h2E1E: out_word = 8'hD5;
		16'h2E1F: out_word = 8'hD9;
		16'h2E20: out_word = 8'hD1;
		16'h2E21: out_word = 8'hD9;
		16'h2E22: out_word = 8'h18;
		16'h2E23: out_word = 8'h57;
		16'h2E24: out_word = 8'hEF;
		16'h2E25: out_word = 8'hE2;
		16'h2E26: out_word = 8'h38;
		16'h2E27: out_word = 8'h7E;
		16'h2E28: out_word = 8'hD6;
		16'h2E29: out_word = 8'h7E;
		16'h2E2A: out_word = 8'hCD;
		16'h2E2B: out_word = 8'hC1;
		16'h2E2C: out_word = 8'h2D;
		16'h2E2D: out_word = 8'h57;
		16'h2E2E: out_word = 8'h3A;
		16'h2E2F: out_word = 8'hAC;
		16'h2E30: out_word = 8'h5C;
		16'h2E31: out_word = 8'h92;
		16'h2E32: out_word = 8'h32;
		16'h2E33: out_word = 8'hAC;
		16'h2E34: out_word = 8'h5C;
		16'h2E35: out_word = 8'h7A;
		16'h2E36: out_word = 8'hCD;
		16'h2E37: out_word = 8'h4F;
		16'h2E38: out_word = 8'h2D;
		16'h2E39: out_word = 8'hEF;
		16'h2E3A: out_word = 8'h31;
		16'h2E3B: out_word = 8'h27;
		16'h2E3C: out_word = 8'hC1;
		16'h2E3D: out_word = 8'h03;
		16'h2E3E: out_word = 8'hE1;
		16'h2E3F: out_word = 8'h38;
		16'h2E40: out_word = 8'hCD;
		16'h2E41: out_word = 8'hD5;
		16'h2E42: out_word = 8'h2D;
		16'h2E43: out_word = 8'hE5;
		16'h2E44: out_word = 8'h32;
		16'h2E45: out_word = 8'hA1;
		16'h2E46: out_word = 8'h5C;
		16'h2E47: out_word = 8'h3D;
		16'h2E48: out_word = 8'h17;
		16'h2E49: out_word = 8'h9F;
		16'h2E4A: out_word = 8'h3C;
		16'h2E4B: out_word = 8'h21;
		16'h2E4C: out_word = 8'hAB;
		16'h2E4D: out_word = 8'h5C;
		16'h2E4E: out_word = 8'h77;
		16'h2E4F: out_word = 8'h23;
		16'h2E50: out_word = 8'h86;
		16'h2E51: out_word = 8'h77;
		16'h2E52: out_word = 8'hE1;
		16'h2E53: out_word = 8'hC3;
		16'h2E54: out_word = 8'hCF;
		16'h2E55: out_word = 8'h2E;
		16'h2E56: out_word = 8'hD6;
		16'h2E57: out_word = 8'h80;
		16'h2E58: out_word = 8'hFE;
		16'h2E59: out_word = 8'h1C;
		16'h2E5A: out_word = 8'h38;
		16'h2E5B: out_word = 8'h13;
		16'h2E5C: out_word = 8'hCD;
		16'h2E5D: out_word = 8'hC1;
		16'h2E5E: out_word = 8'h2D;
		16'h2E5F: out_word = 8'hD6;
		16'h2E60: out_word = 8'h07;
		16'h2E61: out_word = 8'h47;
		16'h2E62: out_word = 8'h21;
		16'h2E63: out_word = 8'hAC;
		16'h2E64: out_word = 8'h5C;
		16'h2E65: out_word = 8'h86;
		16'h2E66: out_word = 8'h77;
		16'h2E67: out_word = 8'h78;
		16'h2E68: out_word = 8'hED;
		16'h2E69: out_word = 8'h44;
		16'h2E6A: out_word = 8'hCD;
		16'h2E6B: out_word = 8'h4F;
		16'h2E6C: out_word = 8'h2D;
		16'h2E6D: out_word = 8'h18;
		16'h2E6E: out_word = 8'h92;
		16'h2E6F: out_word = 8'hEB;
		16'h2E70: out_word = 8'hCD;
		16'h2E71: out_word = 8'hBA;
		16'h2E72: out_word = 8'h2F;
		16'h2E73: out_word = 8'hD9;
		16'h2E74: out_word = 8'hCB;
		16'h2E75: out_word = 8'hFA;
		16'h2E76: out_word = 8'h7D;
		16'h2E77: out_word = 8'hD9;
		16'h2E78: out_word = 8'hD6;
		16'h2E79: out_word = 8'h80;
		16'h2E7A: out_word = 8'h47;
		16'h2E7B: out_word = 8'hCB;
		16'h2E7C: out_word = 8'h23;
		16'h2E7D: out_word = 8'hCB;
		16'h2E7E: out_word = 8'h12;
		16'h2E7F: out_word = 8'hD9;
		16'h2E80: out_word = 8'hCB;
		16'h2E81: out_word = 8'h13;
		16'h2E82: out_word = 8'hCB;
		16'h2E83: out_word = 8'h12;
		16'h2E84: out_word = 8'hD9;
		16'h2E85: out_word = 8'h21;
		16'h2E86: out_word = 8'hAA;
		16'h2E87: out_word = 8'h5C;
		16'h2E88: out_word = 8'h0E;
		16'h2E89: out_word = 8'h05;
		16'h2E8A: out_word = 8'h7E;
		16'h2E8B: out_word = 8'h8F;
		16'h2E8C: out_word = 8'h27;
		16'h2E8D: out_word = 8'h77;
		16'h2E8E: out_word = 8'h2B;
		16'h2E8F: out_word = 8'h0D;
		16'h2E90: out_word = 8'h20;
		16'h2E91: out_word = 8'hF8;
		16'h2E92: out_word = 8'h10;
		16'h2E93: out_word = 8'hE7;
		16'h2E94: out_word = 8'hAF;
		16'h2E95: out_word = 8'h21;
		16'h2E96: out_word = 8'hA6;
		16'h2E97: out_word = 8'h5C;
		16'h2E98: out_word = 8'h11;
		16'h2E99: out_word = 8'hA1;
		16'h2E9A: out_word = 8'h5C;
		16'h2E9B: out_word = 8'h06;
		16'h2E9C: out_word = 8'h09;
		16'h2E9D: out_word = 8'hED;
		16'h2E9E: out_word = 8'h6F;
		16'h2E9F: out_word = 8'h0E;
		16'h2EA0: out_word = 8'hFF;
		16'h2EA1: out_word = 8'hED;
		16'h2EA2: out_word = 8'h6F;
		16'h2EA3: out_word = 8'h20;
		16'h2EA4: out_word = 8'h04;
		16'h2EA5: out_word = 8'h0D;
		16'h2EA6: out_word = 8'h0C;
		16'h2EA7: out_word = 8'h20;
		16'h2EA8: out_word = 8'h0A;
		16'h2EA9: out_word = 8'h12;
		16'h2EAA: out_word = 8'h13;
		16'h2EAB: out_word = 8'hFD;
		16'h2EAC: out_word = 8'h34;
		16'h2EAD: out_word = 8'h71;
		16'h2EAE: out_word = 8'hFD;
		16'h2EAF: out_word = 8'h34;
		16'h2EB0: out_word = 8'h72;
		16'h2EB1: out_word = 8'h0E;
		16'h2EB2: out_word = 8'h00;
		16'h2EB3: out_word = 8'hCB;
		16'h2EB4: out_word = 8'h40;
		16'h2EB5: out_word = 8'h28;
		16'h2EB6: out_word = 8'h01;
		16'h2EB7: out_word = 8'h23;
		16'h2EB8: out_word = 8'h10;
		16'h2EB9: out_word = 8'hE7;
		16'h2EBA: out_word = 8'h3A;
		16'h2EBB: out_word = 8'hAB;
		16'h2EBC: out_word = 8'h5C;
		16'h2EBD: out_word = 8'hD6;
		16'h2EBE: out_word = 8'h09;
		16'h2EBF: out_word = 8'h38;
		16'h2EC0: out_word = 8'h0A;
		16'h2EC1: out_word = 8'hFD;
		16'h2EC2: out_word = 8'h35;
		16'h2EC3: out_word = 8'h71;
		16'h2EC4: out_word = 8'h3E;
		16'h2EC5: out_word = 8'h04;
		16'h2EC6: out_word = 8'hFD;
		16'h2EC7: out_word = 8'hBE;
		16'h2EC8: out_word = 8'h6F;
		16'h2EC9: out_word = 8'h18;
		16'h2ECA: out_word = 8'h41;
		16'h2ECB: out_word = 8'hEF;
		16'h2ECC: out_word = 8'h02;
		16'h2ECD: out_word = 8'hE2;
		16'h2ECE: out_word = 8'h38;
		16'h2ECF: out_word = 8'hEB;
		16'h2ED0: out_word = 8'hCD;
		16'h2ED1: out_word = 8'hBA;
		16'h2ED2: out_word = 8'h2F;
		16'h2ED3: out_word = 8'hD9;
		16'h2ED4: out_word = 8'h3E;
		16'h2ED5: out_word = 8'h80;
		16'h2ED6: out_word = 8'h95;
		16'h2ED7: out_word = 8'h2E;
		16'h2ED8: out_word = 8'h00;
		16'h2ED9: out_word = 8'hCB;
		16'h2EDA: out_word = 8'hFA;
		16'h2EDB: out_word = 8'hD9;
		16'h2EDC: out_word = 8'hCD;
		16'h2EDD: out_word = 8'hDD;
		16'h2EDE: out_word = 8'h2F;
		16'h2EDF: out_word = 8'hFD;
		16'h2EE0: out_word = 8'h7E;
		16'h2EE1: out_word = 8'h71;
		16'h2EE2: out_word = 8'hFE;
		16'h2EE3: out_word = 8'h08;
		16'h2EE4: out_word = 8'h38;
		16'h2EE5: out_word = 8'h06;
		16'h2EE6: out_word = 8'hD9;
		16'h2EE7: out_word = 8'hCB;
		16'h2EE8: out_word = 8'h12;
		16'h2EE9: out_word = 8'hD9;
		16'h2EEA: out_word = 8'h18;
		16'h2EEB: out_word = 8'h20;
		16'h2EEC: out_word = 8'h01;
		16'h2EED: out_word = 8'h00;
		16'h2EEE: out_word = 8'h02;
		16'h2EEF: out_word = 8'h7B;
		16'h2EF0: out_word = 8'hCD;
		16'h2EF1: out_word = 8'h8B;
		16'h2EF2: out_word = 8'h2F;
		16'h2EF3: out_word = 8'h5F;
		16'h2EF4: out_word = 8'h7A;
		16'h2EF5: out_word = 8'hCD;
		16'h2EF6: out_word = 8'h8B;
		16'h2EF7: out_word = 8'h2F;
		16'h2EF8: out_word = 8'h57;
		16'h2EF9: out_word = 8'hC5;
		16'h2EFA: out_word = 8'hD9;
		16'h2EFB: out_word = 8'hC1;
		16'h2EFC: out_word = 8'h10;
		16'h2EFD: out_word = 8'hF1;
		16'h2EFE: out_word = 8'h21;
		16'h2EFF: out_word = 8'hA1;
		16'h2F00: out_word = 8'h5C;
		16'h2F01: out_word = 8'h79;
		16'h2F02: out_word = 8'hFD;
		16'h2F03: out_word = 8'h4E;
		16'h2F04: out_word = 8'h71;
		16'h2F05: out_word = 8'h09;
		16'h2F06: out_word = 8'h77;
		16'h2F07: out_word = 8'hFD;
		16'h2F08: out_word = 8'h34;
		16'h2F09: out_word = 8'h71;
		16'h2F0A: out_word = 8'h18;
		16'h2F0B: out_word = 8'hD3;
		16'h2F0C: out_word = 8'hF5;
		16'h2F0D: out_word = 8'h21;
		16'h2F0E: out_word = 8'hA1;
		16'h2F0F: out_word = 8'h5C;
		16'h2F10: out_word = 8'hFD;
		16'h2F11: out_word = 8'h4E;
		16'h2F12: out_word = 8'h71;
		16'h2F13: out_word = 8'h06;
		16'h2F14: out_word = 8'h00;
		16'h2F15: out_word = 8'h09;
		16'h2F16: out_word = 8'h41;
		16'h2F17: out_word = 8'hF1;
		16'h2F18: out_word = 8'h2B;
		16'h2F19: out_word = 8'h7E;
		16'h2F1A: out_word = 8'hCE;
		16'h2F1B: out_word = 8'h00;
		16'h2F1C: out_word = 8'h77;
		16'h2F1D: out_word = 8'hA7;
		16'h2F1E: out_word = 8'h28;
		16'h2F1F: out_word = 8'h05;
		16'h2F20: out_word = 8'hFE;
		16'h2F21: out_word = 8'h0A;
		16'h2F22: out_word = 8'h3F;
		16'h2F23: out_word = 8'h30;
		16'h2F24: out_word = 8'h08;
		16'h2F25: out_word = 8'h10;
		16'h2F26: out_word = 8'hF1;
		16'h2F27: out_word = 8'h36;
		16'h2F28: out_word = 8'h01;
		16'h2F29: out_word = 8'h04;
		16'h2F2A: out_word = 8'hFD;
		16'h2F2B: out_word = 8'h34;
		16'h2F2C: out_word = 8'h72;
		16'h2F2D: out_word = 8'hFD;
		16'h2F2E: out_word = 8'h70;
		16'h2F2F: out_word = 8'h71;
		16'h2F30: out_word = 8'hEF;
		16'h2F31: out_word = 8'h02;
		16'h2F32: out_word = 8'h38;
		16'h2F33: out_word = 8'hD9;
		16'h2F34: out_word = 8'hE1;
		16'h2F35: out_word = 8'hD9;
		16'h2F36: out_word = 8'hED;
		16'h2F37: out_word = 8'h4B;
		16'h2F38: out_word = 8'hAB;
		16'h2F39: out_word = 8'h5C;
		16'h2F3A: out_word = 8'h21;
		16'h2F3B: out_word = 8'hA1;
		16'h2F3C: out_word = 8'h5C;
		16'h2F3D: out_word = 8'h78;
		16'h2F3E: out_word = 8'hFE;
		16'h2F3F: out_word = 8'h09;
		16'h2F40: out_word = 8'h38;
		16'h2F41: out_word = 8'h04;
		16'h2F42: out_word = 8'hFE;
		16'h2F43: out_word = 8'hFC;
		16'h2F44: out_word = 8'h38;
		16'h2F45: out_word = 8'h26;
		16'h2F46: out_word = 8'hA7;
		16'h2F47: out_word = 8'hCC;
		16'h2F48: out_word = 8'hEF;
		16'h2F49: out_word = 8'h15;
		16'h2F4A: out_word = 8'hAF;
		16'h2F4B: out_word = 8'h90;
		16'h2F4C: out_word = 8'hFA;
		16'h2F4D: out_word = 8'h52;
		16'h2F4E: out_word = 8'h2F;
		16'h2F4F: out_word = 8'h47;
		16'h2F50: out_word = 8'h18;
		16'h2F51: out_word = 8'h0C;
		16'h2F52: out_word = 8'h79;
		16'h2F53: out_word = 8'hA7;
		16'h2F54: out_word = 8'h28;
		16'h2F55: out_word = 8'h03;
		16'h2F56: out_word = 8'h7E;
		16'h2F57: out_word = 8'h23;
		16'h2F58: out_word = 8'h0D;
		16'h2F59: out_word = 8'hCD;
		16'h2F5A: out_word = 8'hEF;
		16'h2F5B: out_word = 8'h15;
		16'h2F5C: out_word = 8'h10;
		16'h2F5D: out_word = 8'hF4;
		16'h2F5E: out_word = 8'h79;
		16'h2F5F: out_word = 8'hA7;
		16'h2F60: out_word = 8'hC8;
		16'h2F61: out_word = 8'h04;
		16'h2F62: out_word = 8'h3E;
		16'h2F63: out_word = 8'h2E;
		16'h2F64: out_word = 8'hD7;
		16'h2F65: out_word = 8'h3E;
		16'h2F66: out_word = 8'h30;
		16'h2F67: out_word = 8'h10;
		16'h2F68: out_word = 8'hFB;
		16'h2F69: out_word = 8'h41;
		16'h2F6A: out_word = 8'h18;
		16'h2F6B: out_word = 8'hE6;
		16'h2F6C: out_word = 8'h50;
		16'h2F6D: out_word = 8'h15;
		16'h2F6E: out_word = 8'h06;
		16'h2F6F: out_word = 8'h01;
		16'h2F70: out_word = 8'hCD;
		16'h2F71: out_word = 8'h4A;
		16'h2F72: out_word = 8'h2F;
		16'h2F73: out_word = 8'h3E;
		16'h2F74: out_word = 8'h45;
		16'h2F75: out_word = 8'hD7;
		16'h2F76: out_word = 8'h4A;
		16'h2F77: out_word = 8'h79;
		16'h2F78: out_word = 8'hA7;
		16'h2F79: out_word = 8'hF2;
		16'h2F7A: out_word = 8'h83;
		16'h2F7B: out_word = 8'h2F;
		16'h2F7C: out_word = 8'hED;
		16'h2F7D: out_word = 8'h44;
		16'h2F7E: out_word = 8'h4F;
		16'h2F7F: out_word = 8'h3E;
		16'h2F80: out_word = 8'h2D;
		16'h2F81: out_word = 8'h18;
		16'h2F82: out_word = 8'h02;
		16'h2F83: out_word = 8'h3E;
		16'h2F84: out_word = 8'h2B;
		16'h2F85: out_word = 8'hD7;
		16'h2F86: out_word = 8'h06;
		16'h2F87: out_word = 8'h00;
		16'h2F88: out_word = 8'hC3;
		16'h2F89: out_word = 8'h1B;
		16'h2F8A: out_word = 8'h1A;
		16'h2F8B: out_word = 8'hD5;
		16'h2F8C: out_word = 8'h6F;
		16'h2F8D: out_word = 8'h26;
		16'h2F8E: out_word = 8'h00;
		16'h2F8F: out_word = 8'h5D;
		16'h2F90: out_word = 8'h54;
		16'h2F91: out_word = 8'h29;
		16'h2F92: out_word = 8'h29;
		16'h2F93: out_word = 8'h19;
		16'h2F94: out_word = 8'h29;
		16'h2F95: out_word = 8'h59;
		16'h2F96: out_word = 8'h19;
		16'h2F97: out_word = 8'h4C;
		16'h2F98: out_word = 8'h7D;
		16'h2F99: out_word = 8'hD1;
		16'h2F9A: out_word = 8'hC9;
		16'h2F9B: out_word = 8'h7E;
		16'h2F9C: out_word = 8'h36;
		16'h2F9D: out_word = 8'h00;
		16'h2F9E: out_word = 8'hA7;
		16'h2F9F: out_word = 8'hC8;
		16'h2FA0: out_word = 8'h23;
		16'h2FA1: out_word = 8'hCB;
		16'h2FA2: out_word = 8'h7E;
		16'h2FA3: out_word = 8'hCB;
		16'h2FA4: out_word = 8'hFE;
		16'h2FA5: out_word = 8'h2B;
		16'h2FA6: out_word = 8'hC8;
		16'h2FA7: out_word = 8'hC5;
		16'h2FA8: out_word = 8'h01;
		16'h2FA9: out_word = 8'h05;
		16'h2FAA: out_word = 8'h00;
		16'h2FAB: out_word = 8'h09;
		16'h2FAC: out_word = 8'h41;
		16'h2FAD: out_word = 8'h4F;
		16'h2FAE: out_word = 8'h37;
		16'h2FAF: out_word = 8'h2B;
		16'h2FB0: out_word = 8'h7E;
		16'h2FB1: out_word = 8'h2F;
		16'h2FB2: out_word = 8'hCE;
		16'h2FB3: out_word = 8'h00;
		16'h2FB4: out_word = 8'h77;
		16'h2FB5: out_word = 8'h10;
		16'h2FB6: out_word = 8'hF8;
		16'h2FB7: out_word = 8'h79;
		16'h2FB8: out_word = 8'hC1;
		16'h2FB9: out_word = 8'hC9;
		16'h2FBA: out_word = 8'hE5;
		16'h2FBB: out_word = 8'hF5;
		16'h2FBC: out_word = 8'h4E;
		16'h2FBD: out_word = 8'h23;
		16'h2FBE: out_word = 8'h46;
		16'h2FBF: out_word = 8'h77;
		16'h2FC0: out_word = 8'h23;
		16'h2FC1: out_word = 8'h79;
		16'h2FC2: out_word = 8'h4E;
		16'h2FC3: out_word = 8'hC5;
		16'h2FC4: out_word = 8'h23;
		16'h2FC5: out_word = 8'h4E;
		16'h2FC6: out_word = 8'h23;
		16'h2FC7: out_word = 8'h46;
		16'h2FC8: out_word = 8'hEB;
		16'h2FC9: out_word = 8'h57;
		16'h2FCA: out_word = 8'h5E;
		16'h2FCB: out_word = 8'hD5;
		16'h2FCC: out_word = 8'h23;
		16'h2FCD: out_word = 8'h56;
		16'h2FCE: out_word = 8'h23;
		16'h2FCF: out_word = 8'h5E;
		16'h2FD0: out_word = 8'hD5;
		16'h2FD1: out_word = 8'hD9;
		16'h2FD2: out_word = 8'hD1;
		16'h2FD3: out_word = 8'hE1;
		16'h2FD4: out_word = 8'hC1;
		16'h2FD5: out_word = 8'hD9;
		16'h2FD6: out_word = 8'h23;
		16'h2FD7: out_word = 8'h56;
		16'h2FD8: out_word = 8'h23;
		16'h2FD9: out_word = 8'h5E;
		16'h2FDA: out_word = 8'hF1;
		16'h2FDB: out_word = 8'hE1;
		16'h2FDC: out_word = 8'hC9;
		16'h2FDD: out_word = 8'hA7;
		16'h2FDE: out_word = 8'hC8;
		16'h2FDF: out_word = 8'hFE;
		16'h2FE0: out_word = 8'h21;
		16'h2FE1: out_word = 8'h30;
		16'h2FE2: out_word = 8'h16;
		16'h2FE3: out_word = 8'hC5;
		16'h2FE4: out_word = 8'h47;
		16'h2FE5: out_word = 8'hD9;
		16'h2FE6: out_word = 8'hCB;
		16'h2FE7: out_word = 8'h2D;
		16'h2FE8: out_word = 8'hCB;
		16'h2FE9: out_word = 8'h1A;
		16'h2FEA: out_word = 8'hCB;
		16'h2FEB: out_word = 8'h1B;
		16'h2FEC: out_word = 8'hD9;
		16'h2FED: out_word = 8'hCB;
		16'h2FEE: out_word = 8'h1A;
		16'h2FEF: out_word = 8'hCB;
		16'h2FF0: out_word = 8'h1B;
		16'h2FF1: out_word = 8'h10;
		16'h2FF2: out_word = 8'hF2;
		16'h2FF3: out_word = 8'hC1;
		16'h2FF4: out_word = 8'hD0;
		16'h2FF5: out_word = 8'hCD;
		16'h2FF6: out_word = 8'h04;
		16'h2FF7: out_word = 8'h30;
		16'h2FF8: out_word = 8'hC0;
		16'h2FF9: out_word = 8'hD9;
		16'h2FFA: out_word = 8'hAF;
		16'h2FFB: out_word = 8'h2E;
		16'h2FFC: out_word = 8'h00;
		16'h2FFD: out_word = 8'h57;
		16'h2FFE: out_word = 8'h5D;
		16'h2FFF: out_word = 8'hD9;
		16'h3000: out_word = 8'h11;
		16'h3001: out_word = 8'h00;
		16'h3002: out_word = 8'h00;
		16'h3003: out_word = 8'hC9;
		16'h3004: out_word = 8'h1C;
		16'h3005: out_word = 8'hC0;
		16'h3006: out_word = 8'h14;
		16'h3007: out_word = 8'hC0;
		16'h3008: out_word = 8'hD9;
		16'h3009: out_word = 8'h1C;
		16'h300A: out_word = 8'h20;
		16'h300B: out_word = 8'h01;
		16'h300C: out_word = 8'h14;
		16'h300D: out_word = 8'hD9;
		16'h300E: out_word = 8'hC9;
		16'h300F: out_word = 8'hEB;
		16'h3010: out_word = 8'hCD;
		16'h3011: out_word = 8'h6E;
		16'h3012: out_word = 8'h34;
		16'h3013: out_word = 8'hEB;
		16'h3014: out_word = 8'h1A;
		16'h3015: out_word = 8'hB6;
		16'h3016: out_word = 8'h20;
		16'h3017: out_word = 8'h26;
		16'h3018: out_word = 8'hD5;
		16'h3019: out_word = 8'h23;
		16'h301A: out_word = 8'hE5;
		16'h301B: out_word = 8'h23;
		16'h301C: out_word = 8'h5E;
		16'h301D: out_word = 8'h23;
		16'h301E: out_word = 8'h56;
		16'h301F: out_word = 8'h23;
		16'h3020: out_word = 8'h23;
		16'h3021: out_word = 8'h23;
		16'h3022: out_word = 8'h7E;
		16'h3023: out_word = 8'h23;
		16'h3024: out_word = 8'h4E;
		16'h3025: out_word = 8'h23;
		16'h3026: out_word = 8'h46;
		16'h3027: out_word = 8'hE1;
		16'h3028: out_word = 8'hEB;
		16'h3029: out_word = 8'h09;
		16'h302A: out_word = 8'hEB;
		16'h302B: out_word = 8'h8E;
		16'h302C: out_word = 8'h0F;
		16'h302D: out_word = 8'hCE;
		16'h302E: out_word = 8'h00;
		16'h302F: out_word = 8'h20;
		16'h3030: out_word = 8'h0B;
		16'h3031: out_word = 8'h9F;
		16'h3032: out_word = 8'h77;
		16'h3033: out_word = 8'h23;
		16'h3034: out_word = 8'h73;
		16'h3035: out_word = 8'h23;
		16'h3036: out_word = 8'h72;
		16'h3037: out_word = 8'h2B;
		16'h3038: out_word = 8'h2B;
		16'h3039: out_word = 8'h2B;
		16'h303A: out_word = 8'hD1;
		16'h303B: out_word = 8'hC9;
		16'h303C: out_word = 8'h2B;
		16'h303D: out_word = 8'hD1;
		16'h303E: out_word = 8'hCD;
		16'h303F: out_word = 8'h93;
		16'h3040: out_word = 8'h32;
		16'h3041: out_word = 8'hD9;
		16'h3042: out_word = 8'hE5;
		16'h3043: out_word = 8'hD9;
		16'h3044: out_word = 8'hD5;
		16'h3045: out_word = 8'hE5;
		16'h3046: out_word = 8'hCD;
		16'h3047: out_word = 8'h9B;
		16'h3048: out_word = 8'h2F;
		16'h3049: out_word = 8'h47;
		16'h304A: out_word = 8'hEB;
		16'h304B: out_word = 8'hCD;
		16'h304C: out_word = 8'h9B;
		16'h304D: out_word = 8'h2F;
		16'h304E: out_word = 8'h4F;
		16'h304F: out_word = 8'hB8;
		16'h3050: out_word = 8'h30;
		16'h3051: out_word = 8'h03;
		16'h3052: out_word = 8'h78;
		16'h3053: out_word = 8'h41;
		16'h3054: out_word = 8'hEB;
		16'h3055: out_word = 8'hF5;
		16'h3056: out_word = 8'h90;
		16'h3057: out_word = 8'hCD;
		16'h3058: out_word = 8'hBA;
		16'h3059: out_word = 8'h2F;
		16'h305A: out_word = 8'hCD;
		16'h305B: out_word = 8'hDD;
		16'h305C: out_word = 8'h2F;
		16'h305D: out_word = 8'hF1;
		16'h305E: out_word = 8'hE1;
		16'h305F: out_word = 8'h77;
		16'h3060: out_word = 8'hE5;
		16'h3061: out_word = 8'h68;
		16'h3062: out_word = 8'h61;
		16'h3063: out_word = 8'h19;
		16'h3064: out_word = 8'hD9;
		16'h3065: out_word = 8'hEB;
		16'h3066: out_word = 8'hED;
		16'h3067: out_word = 8'h4A;
		16'h3068: out_word = 8'hEB;
		16'h3069: out_word = 8'h7C;
		16'h306A: out_word = 8'h8D;
		16'h306B: out_word = 8'h6F;
		16'h306C: out_word = 8'h1F;
		16'h306D: out_word = 8'hAD;
		16'h306E: out_word = 8'hD9;
		16'h306F: out_word = 8'hEB;
		16'h3070: out_word = 8'hE1;
		16'h3071: out_word = 8'h1F;
		16'h3072: out_word = 8'h30;
		16'h3073: out_word = 8'h08;
		16'h3074: out_word = 8'h3E;
		16'h3075: out_word = 8'h01;
		16'h3076: out_word = 8'hCD;
		16'h3077: out_word = 8'hDD;
		16'h3078: out_word = 8'h2F;
		16'h3079: out_word = 8'h34;
		16'h307A: out_word = 8'h28;
		16'h307B: out_word = 8'h23;
		16'h307C: out_word = 8'hD9;
		16'h307D: out_word = 8'h7D;
		16'h307E: out_word = 8'hE6;
		16'h307F: out_word = 8'h80;
		16'h3080: out_word = 8'hD9;
		16'h3081: out_word = 8'h23;
		16'h3082: out_word = 8'h77;
		16'h3083: out_word = 8'h2B;
		16'h3084: out_word = 8'h28;
		16'h3085: out_word = 8'h1F;
		16'h3086: out_word = 8'h7B;
		16'h3087: out_word = 8'hED;
		16'h3088: out_word = 8'h44;
		16'h3089: out_word = 8'h3F;
		16'h308A: out_word = 8'h5F;
		16'h308B: out_word = 8'h7A;
		16'h308C: out_word = 8'h2F;
		16'h308D: out_word = 8'hCE;
		16'h308E: out_word = 8'h00;
		16'h308F: out_word = 8'h57;
		16'h3090: out_word = 8'hD9;
		16'h3091: out_word = 8'h7B;
		16'h3092: out_word = 8'h2F;
		16'h3093: out_word = 8'hCE;
		16'h3094: out_word = 8'h00;
		16'h3095: out_word = 8'h5F;
		16'h3096: out_word = 8'h7A;
		16'h3097: out_word = 8'h2F;
		16'h3098: out_word = 8'hCE;
		16'h3099: out_word = 8'h00;
		16'h309A: out_word = 8'h30;
		16'h309B: out_word = 8'h07;
		16'h309C: out_word = 8'h1F;
		16'h309D: out_word = 8'hD9;
		16'h309E: out_word = 8'h34;
		16'h309F: out_word = 8'hCA;
		16'h30A0: out_word = 8'hAD;
		16'h30A1: out_word = 8'h31;
		16'h30A2: out_word = 8'hD9;
		16'h30A3: out_word = 8'h57;
		16'h30A4: out_word = 8'hD9;
		16'h30A5: out_word = 8'hAF;
		16'h30A6: out_word = 8'hC3;
		16'h30A7: out_word = 8'h55;
		16'h30A8: out_word = 8'h31;
		16'h30A9: out_word = 8'hC5;
		16'h30AA: out_word = 8'h06;
		16'h30AB: out_word = 8'h10;
		16'h30AC: out_word = 8'h7C;
		16'h30AD: out_word = 8'h4D;
		16'h30AE: out_word = 8'h21;
		16'h30AF: out_word = 8'h00;
		16'h30B0: out_word = 8'h00;
		16'h30B1: out_word = 8'h29;
		16'h30B2: out_word = 8'h38;
		16'h30B3: out_word = 8'h0A;
		16'h30B4: out_word = 8'hCB;
		16'h30B5: out_word = 8'h11;
		16'h30B6: out_word = 8'h17;
		16'h30B7: out_word = 8'h30;
		16'h30B8: out_word = 8'h03;
		16'h30B9: out_word = 8'h19;
		16'h30BA: out_word = 8'h38;
		16'h30BB: out_word = 8'h02;
		16'h30BC: out_word = 8'h10;
		16'h30BD: out_word = 8'hF3;
		16'h30BE: out_word = 8'hC1;
		16'h30BF: out_word = 8'hC9;
		16'h30C0: out_word = 8'hCD;
		16'h30C1: out_word = 8'hE9;
		16'h30C2: out_word = 8'h34;
		16'h30C3: out_word = 8'hD8;
		16'h30C4: out_word = 8'h23;
		16'h30C5: out_word = 8'hAE;
		16'h30C6: out_word = 8'hCB;
		16'h30C7: out_word = 8'hFE;
		16'h30C8: out_word = 8'h2B;
		16'h30C9: out_word = 8'hC9;
		16'h30CA: out_word = 8'h1A;
		16'h30CB: out_word = 8'hB6;
		16'h30CC: out_word = 8'h20;
		16'h30CD: out_word = 8'h22;
		16'h30CE: out_word = 8'hD5;
		16'h30CF: out_word = 8'hE5;
		16'h30D0: out_word = 8'hD5;
		16'h30D1: out_word = 8'hCD;
		16'h30D2: out_word = 8'h7F;
		16'h30D3: out_word = 8'h2D;
		16'h30D4: out_word = 8'hEB;
		16'h30D5: out_word = 8'hE3;
		16'h30D6: out_word = 8'h41;
		16'h30D7: out_word = 8'hCD;
		16'h30D8: out_word = 8'h7F;
		16'h30D9: out_word = 8'h2D;
		16'h30DA: out_word = 8'h78;
		16'h30DB: out_word = 8'hA9;
		16'h30DC: out_word = 8'h4F;
		16'h30DD: out_word = 8'hE1;
		16'h30DE: out_word = 8'hCD;
		16'h30DF: out_word = 8'hA9;
		16'h30E0: out_word = 8'h30;
		16'h30E1: out_word = 8'hEB;
		16'h30E2: out_word = 8'hE1;
		16'h30E3: out_word = 8'h38;
		16'h30E4: out_word = 8'h0A;
		16'h30E5: out_word = 8'h7A;
		16'h30E6: out_word = 8'hB3;
		16'h30E7: out_word = 8'h20;
		16'h30E8: out_word = 8'h01;
		16'h30E9: out_word = 8'h4F;
		16'h30EA: out_word = 8'hCD;
		16'h30EB: out_word = 8'h8E;
		16'h30EC: out_word = 8'h2D;
		16'h30ED: out_word = 8'hD1;
		16'h30EE: out_word = 8'hC9;
		16'h30EF: out_word = 8'hD1;
		16'h30F0: out_word = 8'hCD;
		16'h30F1: out_word = 8'h93;
		16'h30F2: out_word = 8'h32;
		16'h30F3: out_word = 8'hAF;
		16'h30F4: out_word = 8'hCD;
		16'h30F5: out_word = 8'hC0;
		16'h30F6: out_word = 8'h30;
		16'h30F7: out_word = 8'hD8;
		16'h30F8: out_word = 8'hD9;
		16'h30F9: out_word = 8'hE5;
		16'h30FA: out_word = 8'hD9;
		16'h30FB: out_word = 8'hD5;
		16'h30FC: out_word = 8'hEB;
		16'h30FD: out_word = 8'hCD;
		16'h30FE: out_word = 8'hC0;
		16'h30FF: out_word = 8'h30;
		16'h3100: out_word = 8'hEB;
		16'h3101: out_word = 8'h38;
		16'h3102: out_word = 8'h5A;
		16'h3103: out_word = 8'hE5;
		16'h3104: out_word = 8'hCD;
		16'h3105: out_word = 8'hBA;
		16'h3106: out_word = 8'h2F;
		16'h3107: out_word = 8'h78;
		16'h3108: out_word = 8'hA7;
		16'h3109: out_word = 8'hED;
		16'h310A: out_word = 8'h62;
		16'h310B: out_word = 8'hD9;
		16'h310C: out_word = 8'hE5;
		16'h310D: out_word = 8'hED;
		16'h310E: out_word = 8'h62;
		16'h310F: out_word = 8'hD9;
		16'h3110: out_word = 8'h06;
		16'h3111: out_word = 8'h21;
		16'h3112: out_word = 8'h18;
		16'h3113: out_word = 8'h11;
		16'h3114: out_word = 8'h30;
		16'h3115: out_word = 8'h05;
		16'h3116: out_word = 8'h19;
		16'h3117: out_word = 8'hD9;
		16'h3118: out_word = 8'hED;
		16'h3119: out_word = 8'h5A;
		16'h311A: out_word = 8'hD9;
		16'h311B: out_word = 8'hD9;
		16'h311C: out_word = 8'hCB;
		16'h311D: out_word = 8'h1C;
		16'h311E: out_word = 8'hCB;
		16'h311F: out_word = 8'h1D;
		16'h3120: out_word = 8'hD9;
		16'h3121: out_word = 8'hCB;
		16'h3122: out_word = 8'h1C;
		16'h3123: out_word = 8'hCB;
		16'h3124: out_word = 8'h1D;
		16'h3125: out_word = 8'hD9;
		16'h3126: out_word = 8'hCB;
		16'h3127: out_word = 8'h18;
		16'h3128: out_word = 8'hCB;
		16'h3129: out_word = 8'h19;
		16'h312A: out_word = 8'hD9;
		16'h312B: out_word = 8'hCB;
		16'h312C: out_word = 8'h19;
		16'h312D: out_word = 8'h1F;
		16'h312E: out_word = 8'h10;
		16'h312F: out_word = 8'hE4;
		16'h3130: out_word = 8'hEB;
		16'h3131: out_word = 8'hD9;
		16'h3132: out_word = 8'hEB;
		16'h3133: out_word = 8'hD9;
		16'h3134: out_word = 8'hC1;
		16'h3135: out_word = 8'hE1;
		16'h3136: out_word = 8'h78;
		16'h3137: out_word = 8'h81;
		16'h3138: out_word = 8'h20;
		16'h3139: out_word = 8'h01;
		16'h313A: out_word = 8'hA7;
		16'h313B: out_word = 8'h3D;
		16'h313C: out_word = 8'h3F;
		16'h313D: out_word = 8'h17;
		16'h313E: out_word = 8'h3F;
		16'h313F: out_word = 8'h1F;
		16'h3140: out_word = 8'hF2;
		16'h3141: out_word = 8'h46;
		16'h3142: out_word = 8'h31;
		16'h3143: out_word = 8'h30;
		16'h3144: out_word = 8'h68;
		16'h3145: out_word = 8'hA7;
		16'h3146: out_word = 8'h3C;
		16'h3147: out_word = 8'h20;
		16'h3148: out_word = 8'h08;
		16'h3149: out_word = 8'h38;
		16'h314A: out_word = 8'h06;
		16'h314B: out_word = 8'hD9;
		16'h314C: out_word = 8'hCB;
		16'h314D: out_word = 8'h7A;
		16'h314E: out_word = 8'hD9;
		16'h314F: out_word = 8'h20;
		16'h3150: out_word = 8'h5C;
		16'h3151: out_word = 8'h77;
		16'h3152: out_word = 8'hD9;
		16'h3153: out_word = 8'h78;
		16'h3154: out_word = 8'hD9;
		16'h3155: out_word = 8'h30;
		16'h3156: out_word = 8'h15;
		16'h3157: out_word = 8'h7E;
		16'h3158: out_word = 8'hA7;
		16'h3159: out_word = 8'h3E;
		16'h315A: out_word = 8'h80;
		16'h315B: out_word = 8'h28;
		16'h315C: out_word = 8'h01;
		16'h315D: out_word = 8'hAF;
		16'h315E: out_word = 8'hD9;
		16'h315F: out_word = 8'hA2;
		16'h3160: out_word = 8'hCD;
		16'h3161: out_word = 8'hFB;
		16'h3162: out_word = 8'h2F;
		16'h3163: out_word = 8'h07;
		16'h3164: out_word = 8'h77;
		16'h3165: out_word = 8'h38;
		16'h3166: out_word = 8'h2E;
		16'h3167: out_word = 8'h23;
		16'h3168: out_word = 8'h77;
		16'h3169: out_word = 8'h2B;
		16'h316A: out_word = 8'h18;
		16'h316B: out_word = 8'h29;
		16'h316C: out_word = 8'h06;
		16'h316D: out_word = 8'h20;
		16'h316E: out_word = 8'hD9;
		16'h316F: out_word = 8'hCB;
		16'h3170: out_word = 8'h7A;
		16'h3171: out_word = 8'hD9;
		16'h3172: out_word = 8'h20;
		16'h3173: out_word = 8'h12;
		16'h3174: out_word = 8'h07;
		16'h3175: out_word = 8'hCB;
		16'h3176: out_word = 8'h13;
		16'h3177: out_word = 8'hCB;
		16'h3178: out_word = 8'h12;
		16'h3179: out_word = 8'hD9;
		16'h317A: out_word = 8'hCB;
		16'h317B: out_word = 8'h13;
		16'h317C: out_word = 8'hCB;
		16'h317D: out_word = 8'h12;
		16'h317E: out_word = 8'hD9;
		16'h317F: out_word = 8'h35;
		16'h3180: out_word = 8'h28;
		16'h3181: out_word = 8'hD7;
		16'h3182: out_word = 8'h10;
		16'h3183: out_word = 8'hEA;
		16'h3184: out_word = 8'h18;
		16'h3185: out_word = 8'hD7;
		16'h3186: out_word = 8'h17;
		16'h3187: out_word = 8'h30;
		16'h3188: out_word = 8'h0C;
		16'h3189: out_word = 8'hCD;
		16'h318A: out_word = 8'h04;
		16'h318B: out_word = 8'h30;
		16'h318C: out_word = 8'h20;
		16'h318D: out_word = 8'h07;
		16'h318E: out_word = 8'hD9;
		16'h318F: out_word = 8'h16;
		16'h3190: out_word = 8'h80;
		16'h3191: out_word = 8'hD9;
		16'h3192: out_word = 8'h34;
		16'h3193: out_word = 8'h28;
		16'h3194: out_word = 8'h18;
		16'h3195: out_word = 8'hE5;
		16'h3196: out_word = 8'h23;
		16'h3197: out_word = 8'hD9;
		16'h3198: out_word = 8'hD5;
		16'h3199: out_word = 8'hD9;
		16'h319A: out_word = 8'hC1;
		16'h319B: out_word = 8'h78;
		16'h319C: out_word = 8'h17;
		16'h319D: out_word = 8'hCB;
		16'h319E: out_word = 8'h16;
		16'h319F: out_word = 8'h1F;
		16'h31A0: out_word = 8'h77;
		16'h31A1: out_word = 8'h23;
		16'h31A2: out_word = 8'h71;
		16'h31A3: out_word = 8'h23;
		16'h31A4: out_word = 8'h72;
		16'h31A5: out_word = 8'h23;
		16'h31A6: out_word = 8'h73;
		16'h31A7: out_word = 8'hE1;
		16'h31A8: out_word = 8'hD1;
		16'h31A9: out_word = 8'hD9;
		16'h31AA: out_word = 8'hE1;
		16'h31AB: out_word = 8'hD9;
		16'h31AC: out_word = 8'hC9;
		16'h31AD: out_word = 8'hCF;
		16'h31AE: out_word = 8'h05;
		16'h31AF: out_word = 8'hCD;
		16'h31B0: out_word = 8'h93;
		16'h31B1: out_word = 8'h32;
		16'h31B2: out_word = 8'hEB;
		16'h31B3: out_word = 8'hAF;
		16'h31B4: out_word = 8'hCD;
		16'h31B5: out_word = 8'hC0;
		16'h31B6: out_word = 8'h30;
		16'h31B7: out_word = 8'h38;
		16'h31B8: out_word = 8'hF4;
		16'h31B9: out_word = 8'hEB;
		16'h31BA: out_word = 8'hCD;
		16'h31BB: out_word = 8'hC0;
		16'h31BC: out_word = 8'h30;
		16'h31BD: out_word = 8'hD8;
		16'h31BE: out_word = 8'hD9;
		16'h31BF: out_word = 8'hE5;
		16'h31C0: out_word = 8'hD9;
		16'h31C1: out_word = 8'hD5;
		16'h31C2: out_word = 8'hE5;
		16'h31C3: out_word = 8'hCD;
		16'h31C4: out_word = 8'hBA;
		16'h31C5: out_word = 8'h2F;
		16'h31C6: out_word = 8'hD9;
		16'h31C7: out_word = 8'hE5;
		16'h31C8: out_word = 8'h60;
		16'h31C9: out_word = 8'h69;
		16'h31CA: out_word = 8'hD9;
		16'h31CB: out_word = 8'h61;
		16'h31CC: out_word = 8'h68;
		16'h31CD: out_word = 8'hAF;
		16'h31CE: out_word = 8'h06;
		16'h31CF: out_word = 8'hDF;
		16'h31D0: out_word = 8'h18;
		16'h31D1: out_word = 8'h10;
		16'h31D2: out_word = 8'h17;
		16'h31D3: out_word = 8'hCB;
		16'h31D4: out_word = 8'h11;
		16'h31D5: out_word = 8'hD9;
		16'h31D6: out_word = 8'hCB;
		16'h31D7: out_word = 8'h11;
		16'h31D8: out_word = 8'hCB;
		16'h31D9: out_word = 8'h10;
		16'h31DA: out_word = 8'hD9;
		16'h31DB: out_word = 8'h29;
		16'h31DC: out_word = 8'hD9;
		16'h31DD: out_word = 8'hED;
		16'h31DE: out_word = 8'h6A;
		16'h31DF: out_word = 8'hD9;
		16'h31E0: out_word = 8'h38;
		16'h31E1: out_word = 8'h10;
		16'h31E2: out_word = 8'hED;
		16'h31E3: out_word = 8'h52;
		16'h31E4: out_word = 8'hD9;
		16'h31E5: out_word = 8'hED;
		16'h31E6: out_word = 8'h52;
		16'h31E7: out_word = 8'hD9;
		16'h31E8: out_word = 8'h30;
		16'h31E9: out_word = 8'h0F;
		16'h31EA: out_word = 8'h19;
		16'h31EB: out_word = 8'hD9;
		16'h31EC: out_word = 8'hED;
		16'h31ED: out_word = 8'h5A;
		16'h31EE: out_word = 8'hD9;
		16'h31EF: out_word = 8'hA7;
		16'h31F0: out_word = 8'h18;
		16'h31F1: out_word = 8'h08;
		16'h31F2: out_word = 8'hA7;
		16'h31F3: out_word = 8'hED;
		16'h31F4: out_word = 8'h52;
		16'h31F5: out_word = 8'hD9;
		16'h31F6: out_word = 8'hED;
		16'h31F7: out_word = 8'h52;
		16'h31F8: out_word = 8'hD9;
		16'h31F9: out_word = 8'h37;
		16'h31FA: out_word = 8'h04;
		16'h31FB: out_word = 8'hFA;
		16'h31FC: out_word = 8'hD2;
		16'h31FD: out_word = 8'h31;
		16'h31FE: out_word = 8'hF5;
		16'h31FF: out_word = 8'h28;
		16'h3200: out_word = 8'hE1;
		16'h3201: out_word = 8'h5F;
		16'h3202: out_word = 8'h51;
		16'h3203: out_word = 8'hD9;
		16'h3204: out_word = 8'h59;
		16'h3205: out_word = 8'h50;
		16'h3206: out_word = 8'hF1;
		16'h3207: out_word = 8'hCB;
		16'h3208: out_word = 8'h18;
		16'h3209: out_word = 8'hF1;
		16'h320A: out_word = 8'hCB;
		16'h320B: out_word = 8'h18;
		16'h320C: out_word = 8'hD9;
		16'h320D: out_word = 8'hC1;
		16'h320E: out_word = 8'hE1;
		16'h320F: out_word = 8'h78;
		16'h3210: out_word = 8'h91;
		16'h3211: out_word = 8'hC3;
		16'h3212: out_word = 8'h3D;
		16'h3213: out_word = 8'h31;
		16'h3214: out_word = 8'h7E;
		16'h3215: out_word = 8'hA7;
		16'h3216: out_word = 8'hC8;
		16'h3217: out_word = 8'hFE;
		16'h3218: out_word = 8'h81;
		16'h3219: out_word = 8'h30;
		16'h321A: out_word = 8'h06;
		16'h321B: out_word = 8'h36;
		16'h321C: out_word = 8'h00;
		16'h321D: out_word = 8'h3E;
		16'h321E: out_word = 8'h20;
		16'h321F: out_word = 8'h18;
		16'h3220: out_word = 8'h51;
		16'h3221: out_word = 8'hFE;
		16'h3222: out_word = 8'h91;
		16'h3223: out_word = 8'h20;
		16'h3224: out_word = 8'h1A;
		16'h3225: out_word = 8'h23;
		16'h3226: out_word = 8'h23;
		16'h3227: out_word = 8'h23;
		16'h3228: out_word = 8'h3E;
		16'h3229: out_word = 8'h80;
		16'h322A: out_word = 8'hA6;
		16'h322B: out_word = 8'h2B;
		16'h322C: out_word = 8'hB6;
		16'h322D: out_word = 8'h2B;
		16'h322E: out_word = 8'h20;
		16'h322F: out_word = 8'h03;
		16'h3230: out_word = 8'h3E;
		16'h3231: out_word = 8'h80;
		16'h3232: out_word = 8'hAE;
		16'h3233: out_word = 8'h2B;
		16'h3234: out_word = 8'h20;
		16'h3235: out_word = 8'h36;
		16'h3236: out_word = 8'h77;
		16'h3237: out_word = 8'h23;
		16'h3238: out_word = 8'h36;
		16'h3239: out_word = 8'hFF;
		16'h323A: out_word = 8'h2B;
		16'h323B: out_word = 8'h3E;
		16'h323C: out_word = 8'h18;
		16'h323D: out_word = 8'h18;
		16'h323E: out_word = 8'h33;
		16'h323F: out_word = 8'h30;
		16'h3240: out_word = 8'h2C;
		16'h3241: out_word = 8'hD5;
		16'h3242: out_word = 8'h2F;
		16'h3243: out_word = 8'hC6;
		16'h3244: out_word = 8'h91;
		16'h3245: out_word = 8'h23;
		16'h3246: out_word = 8'h56;
		16'h3247: out_word = 8'h23;
		16'h3248: out_word = 8'h5E;
		16'h3249: out_word = 8'h2B;
		16'h324A: out_word = 8'h2B;
		16'h324B: out_word = 8'h0E;
		16'h324C: out_word = 8'h00;
		16'h324D: out_word = 8'hCB;
		16'h324E: out_word = 8'h7A;
		16'h324F: out_word = 8'h28;
		16'h3250: out_word = 8'h01;
		16'h3251: out_word = 8'h0D;
		16'h3252: out_word = 8'hCB;
		16'h3253: out_word = 8'hFA;
		16'h3254: out_word = 8'h06;
		16'h3255: out_word = 8'h08;
		16'h3256: out_word = 8'h90;
		16'h3257: out_word = 8'h80;
		16'h3258: out_word = 8'h38;
		16'h3259: out_word = 8'h04;
		16'h325A: out_word = 8'h5A;
		16'h325B: out_word = 8'h16;
		16'h325C: out_word = 8'h00;
		16'h325D: out_word = 8'h90;
		16'h325E: out_word = 8'h28;
		16'h325F: out_word = 8'h07;
		16'h3260: out_word = 8'h47;
		16'h3261: out_word = 8'hCB;
		16'h3262: out_word = 8'h3A;
		16'h3263: out_word = 8'hCB;
		16'h3264: out_word = 8'h1B;
		16'h3265: out_word = 8'h10;
		16'h3266: out_word = 8'hFA;
		16'h3267: out_word = 8'hCD;
		16'h3268: out_word = 8'h8E;
		16'h3269: out_word = 8'h2D;
		16'h326A: out_word = 8'hD1;
		16'h326B: out_word = 8'hC9;
		16'h326C: out_word = 8'h7E;
		16'h326D: out_word = 8'hD6;
		16'h326E: out_word = 8'hA0;
		16'h326F: out_word = 8'hF0;
		16'h3270: out_word = 8'hED;
		16'h3271: out_word = 8'h44;
		16'h3272: out_word = 8'hD5;
		16'h3273: out_word = 8'hEB;
		16'h3274: out_word = 8'h2B;
		16'h3275: out_word = 8'h47;
		16'h3276: out_word = 8'hCB;
		16'h3277: out_word = 8'h38;
		16'h3278: out_word = 8'hCB;
		16'h3279: out_word = 8'h38;
		16'h327A: out_word = 8'hCB;
		16'h327B: out_word = 8'h38;
		16'h327C: out_word = 8'h28;
		16'h327D: out_word = 8'h05;
		16'h327E: out_word = 8'h36;
		16'h327F: out_word = 8'h00;
		16'h3280: out_word = 8'h2B;
		16'h3281: out_word = 8'h10;
		16'h3282: out_word = 8'hFB;
		16'h3283: out_word = 8'hE6;
		16'h3284: out_word = 8'h07;
		16'h3285: out_word = 8'h28;
		16'h3286: out_word = 8'h09;
		16'h3287: out_word = 8'h47;
		16'h3288: out_word = 8'h3E;
		16'h3289: out_word = 8'hFF;
		16'h328A: out_word = 8'hCB;
		16'h328B: out_word = 8'h27;
		16'h328C: out_word = 8'h10;
		16'h328D: out_word = 8'hFC;
		16'h328E: out_word = 8'hA6;
		16'h328F: out_word = 8'h77;
		16'h3290: out_word = 8'hEB;
		16'h3291: out_word = 8'hD1;
		16'h3292: out_word = 8'hC9;
		16'h3293: out_word = 8'hCD;
		16'h3294: out_word = 8'h96;
		16'h3295: out_word = 8'h32;
		16'h3296: out_word = 8'hEB;
		16'h3297: out_word = 8'h7E;
		16'h3298: out_word = 8'hA7;
		16'h3299: out_word = 8'hC0;
		16'h329A: out_word = 8'hD5;
		16'h329B: out_word = 8'hCD;
		16'h329C: out_word = 8'h7F;
		16'h329D: out_word = 8'h2D;
		16'h329E: out_word = 8'hAF;
		16'h329F: out_word = 8'h23;
		16'h32A0: out_word = 8'h77;
		16'h32A1: out_word = 8'h2B;
		16'h32A2: out_word = 8'h77;
		16'h32A3: out_word = 8'h06;
		16'h32A4: out_word = 8'h91;
		16'h32A5: out_word = 8'h7A;
		16'h32A6: out_word = 8'hA7;
		16'h32A7: out_word = 8'h20;
		16'h32A8: out_word = 8'h08;
		16'h32A9: out_word = 8'hB3;
		16'h32AA: out_word = 8'h42;
		16'h32AB: out_word = 8'h28;
		16'h32AC: out_word = 8'h10;
		16'h32AD: out_word = 8'h53;
		16'h32AE: out_word = 8'h58;
		16'h32AF: out_word = 8'h06;
		16'h32B0: out_word = 8'h89;
		16'h32B1: out_word = 8'hEB;
		16'h32B2: out_word = 8'h05;
		16'h32B3: out_word = 8'h29;
		16'h32B4: out_word = 8'h30;
		16'h32B5: out_word = 8'hFC;
		16'h32B6: out_word = 8'hCB;
		16'h32B7: out_word = 8'h09;
		16'h32B8: out_word = 8'hCB;
		16'h32B9: out_word = 8'h1C;
		16'h32BA: out_word = 8'hCB;
		16'h32BB: out_word = 8'h1D;
		16'h32BC: out_word = 8'hEB;
		16'h32BD: out_word = 8'h2B;
		16'h32BE: out_word = 8'h73;
		16'h32BF: out_word = 8'h2B;
		16'h32C0: out_word = 8'h72;
		16'h32C1: out_word = 8'h2B;
		16'h32C2: out_word = 8'h70;
		16'h32C3: out_word = 8'hD1;
		16'h32C4: out_word = 8'hC9;
		16'h32C5: out_word = 8'h00;
		16'h32C6: out_word = 8'hB0;
		16'h32C7: out_word = 8'h00;
		16'h32C8: out_word = 8'h40;
		16'h32C9: out_word = 8'hB0;
		16'h32CA: out_word = 8'h00;
		16'h32CB: out_word = 8'h01;
		16'h32CC: out_word = 8'h30;
		16'h32CD: out_word = 8'h00;
		16'h32CE: out_word = 8'hF1;
		16'h32CF: out_word = 8'h49;
		16'h32D0: out_word = 8'h0F;
		16'h32D1: out_word = 8'hDA;
		16'h32D2: out_word = 8'hA2;
		16'h32D3: out_word = 8'h40;
		16'h32D4: out_word = 8'hB0;
		16'h32D5: out_word = 8'h00;
		16'h32D6: out_word = 8'h0A;
		16'h32D7: out_word = 8'h8F;
		16'h32D8: out_word = 8'h36;
		16'h32D9: out_word = 8'h3C;
		16'h32DA: out_word = 8'h34;
		16'h32DB: out_word = 8'hA1;
		16'h32DC: out_word = 8'h33;
		16'h32DD: out_word = 8'h0F;
		16'h32DE: out_word = 8'h30;
		16'h32DF: out_word = 8'hCA;
		16'h32E0: out_word = 8'h30;
		16'h32E1: out_word = 8'hAF;
		16'h32E2: out_word = 8'h31;
		16'h32E3: out_word = 8'h51;
		16'h32E4: out_word = 8'h38;
		16'h32E5: out_word = 8'h1B;
		16'h32E6: out_word = 8'h35;
		16'h32E7: out_word = 8'h24;
		16'h32E8: out_word = 8'h35;
		16'h32E9: out_word = 8'h3B;
		16'h32EA: out_word = 8'h35;
		16'h32EB: out_word = 8'h3B;
		16'h32EC: out_word = 8'h35;
		16'h32ED: out_word = 8'h3B;
		16'h32EE: out_word = 8'h35;
		16'h32EF: out_word = 8'h3B;
		16'h32F0: out_word = 8'h35;
		16'h32F1: out_word = 8'h3B;
		16'h32F2: out_word = 8'h35;
		16'h32F3: out_word = 8'h3B;
		16'h32F4: out_word = 8'h35;
		16'h32F5: out_word = 8'h14;
		16'h32F6: out_word = 8'h30;
		16'h32F7: out_word = 8'h2D;
		16'h32F8: out_word = 8'h35;
		16'h32F9: out_word = 8'h3B;
		16'h32FA: out_word = 8'h35;
		16'h32FB: out_word = 8'h3B;
		16'h32FC: out_word = 8'h35;
		16'h32FD: out_word = 8'h3B;
		16'h32FE: out_word = 8'h35;
		16'h32FF: out_word = 8'h3B;
		16'h3300: out_word = 8'h35;
		16'h3301: out_word = 8'h3B;
		16'h3302: out_word = 8'h35;
		16'h3303: out_word = 8'h3B;
		16'h3304: out_word = 8'h35;
		16'h3305: out_word = 8'h9C;
		16'h3306: out_word = 8'h35;
		16'h3307: out_word = 8'hDE;
		16'h3308: out_word = 8'h35;
		16'h3309: out_word = 8'hBC;
		16'h330A: out_word = 8'h34;
		16'h330B: out_word = 8'h45;
		16'h330C: out_word = 8'h36;
		16'h330D: out_word = 8'h6E;
		16'h330E: out_word = 8'h34;
		16'h330F: out_word = 8'h69;
		16'h3310: out_word = 8'h36;
		16'h3311: out_word = 8'hDE;
		16'h3312: out_word = 8'h35;
		16'h3313: out_word = 8'h74;
		16'h3314: out_word = 8'h36;
		16'h3315: out_word = 8'hB5;
		16'h3316: out_word = 8'h37;
		16'h3317: out_word = 8'hAA;
		16'h3318: out_word = 8'h37;
		16'h3319: out_word = 8'hDA;
		16'h331A: out_word = 8'h37;
		16'h331B: out_word = 8'h33;
		16'h331C: out_word = 8'h38;
		16'h331D: out_word = 8'h43;
		16'h331E: out_word = 8'h38;
		16'h331F: out_word = 8'hE2;
		16'h3320: out_word = 8'h37;
		16'h3321: out_word = 8'h13;
		16'h3322: out_word = 8'h37;
		16'h3323: out_word = 8'hC4;
		16'h3324: out_word = 8'h36;
		16'h3325: out_word = 8'hAF;
		16'h3326: out_word = 8'h36;
		16'h3327: out_word = 8'h4A;
		16'h3328: out_word = 8'h38;
		16'h3329: out_word = 8'h92;
		16'h332A: out_word = 8'h34;
		16'h332B: out_word = 8'h6A;
		16'h332C: out_word = 8'h34;
		16'h332D: out_word = 8'hAC;
		16'h332E: out_word = 8'h34;
		16'h332F: out_word = 8'hA5;
		16'h3330: out_word = 8'h34;
		16'h3331: out_word = 8'hB3;
		16'h3332: out_word = 8'h34;
		16'h3333: out_word = 8'h1F;
		16'h3334: out_word = 8'h36;
		16'h3335: out_word = 8'hC9;
		16'h3336: out_word = 8'h35;
		16'h3337: out_word = 8'h01;
		16'h3338: out_word = 8'h35;
		16'h3339: out_word = 8'hC0;
		16'h333A: out_word = 8'h33;
		16'h333B: out_word = 8'hA0;
		16'h333C: out_word = 8'h36;
		16'h333D: out_word = 8'h86;
		16'h333E: out_word = 8'h36;
		16'h333F: out_word = 8'hC6;
		16'h3340: out_word = 8'h33;
		16'h3341: out_word = 8'h7A;
		16'h3342: out_word = 8'h36;
		16'h3343: out_word = 8'h06;
		16'h3344: out_word = 8'h35;
		16'h3345: out_word = 8'hF9;
		16'h3346: out_word = 8'h34;
		16'h3347: out_word = 8'h9B;
		16'h3348: out_word = 8'h36;
		16'h3349: out_word = 8'h83;
		16'h334A: out_word = 8'h37;
		16'h334B: out_word = 8'h14;
		16'h334C: out_word = 8'h32;
		16'h334D: out_word = 8'hA2;
		16'h334E: out_word = 8'h33;
		16'h334F: out_word = 8'h4F;
		16'h3350: out_word = 8'h2D;
		16'h3351: out_word = 8'h97;
		16'h3352: out_word = 8'h32;
		16'h3353: out_word = 8'h49;
		16'h3354: out_word = 8'h34;
		16'h3355: out_word = 8'h1B;
		16'h3356: out_word = 8'h34;
		16'h3357: out_word = 8'h2D;
		16'h3358: out_word = 8'h34;
		16'h3359: out_word = 8'h0F;
		16'h335A: out_word = 8'h34;
		16'h335B: out_word = 8'hCD;
		16'h335C: out_word = 8'hBF;
		16'h335D: out_word = 8'h35;
		16'h335E: out_word = 8'h78;
		16'h335F: out_word = 8'h32;
		16'h3360: out_word = 8'h67;
		16'h3361: out_word = 8'h5C;
		16'h3362: out_word = 8'hD9;
		16'h3363: out_word = 8'hE3;
		16'h3364: out_word = 8'hD9;
		16'h3365: out_word = 8'hED;
		16'h3366: out_word = 8'h53;
		16'h3367: out_word = 8'h65;
		16'h3368: out_word = 8'h5C;
		16'h3369: out_word = 8'hD9;
		16'h336A: out_word = 8'h7E;
		16'h336B: out_word = 8'h23;
		16'h336C: out_word = 8'hE5;
		16'h336D: out_word = 8'hA7;
		16'h336E: out_word = 8'hF2;
		16'h336F: out_word = 8'h80;
		16'h3370: out_word = 8'h33;
		16'h3371: out_word = 8'h57;
		16'h3372: out_word = 8'hE6;
		16'h3373: out_word = 8'h60;
		16'h3374: out_word = 8'h0F;
		16'h3375: out_word = 8'h0F;
		16'h3376: out_word = 8'h0F;
		16'h3377: out_word = 8'h0F;
		16'h3378: out_word = 8'hC6;
		16'h3379: out_word = 8'h7C;
		16'h337A: out_word = 8'h6F;
		16'h337B: out_word = 8'h7A;
		16'h337C: out_word = 8'hE6;
		16'h337D: out_word = 8'h1F;
		16'h337E: out_word = 8'h18;
		16'h337F: out_word = 8'h0E;
		16'h3380: out_word = 8'hFE;
		16'h3381: out_word = 8'h18;
		16'h3382: out_word = 8'h30;
		16'h3383: out_word = 8'h08;
		16'h3384: out_word = 8'hD9;
		16'h3385: out_word = 8'h01;
		16'h3386: out_word = 8'hFB;
		16'h3387: out_word = 8'hFF;
		16'h3388: out_word = 8'h54;
		16'h3389: out_word = 8'h5D;
		16'h338A: out_word = 8'h09;
		16'h338B: out_word = 8'hD9;
		16'h338C: out_word = 8'h07;
		16'h338D: out_word = 8'h6F;
		16'h338E: out_word = 8'h11;
		16'h338F: out_word = 8'hD7;
		16'h3390: out_word = 8'h32;
		16'h3391: out_word = 8'h26;
		16'h3392: out_word = 8'h00;
		16'h3393: out_word = 8'h19;
		16'h3394: out_word = 8'h5E;
		16'h3395: out_word = 8'h23;
		16'h3396: out_word = 8'h56;
		16'h3397: out_word = 8'h21;
		16'h3398: out_word = 8'h65;
		16'h3399: out_word = 8'h33;
		16'h339A: out_word = 8'hE3;
		16'h339B: out_word = 8'hD5;
		16'h339C: out_word = 8'hD9;
		16'h339D: out_word = 8'hED;
		16'h339E: out_word = 8'h4B;
		16'h339F: out_word = 8'h66;
		16'h33A0: out_word = 8'h5C;
		16'h33A1: out_word = 8'hC9;
		16'h33A2: out_word = 8'hF1;
		16'h33A3: out_word = 8'h3A;
		16'h33A4: out_word = 8'h67;
		16'h33A5: out_word = 8'h5C;
		16'h33A6: out_word = 8'hD9;
		16'h33A7: out_word = 8'h18;
		16'h33A8: out_word = 8'hC3;
		16'h33A9: out_word = 8'hD5;
		16'h33AA: out_word = 8'hE5;
		16'h33AB: out_word = 8'h01;
		16'h33AC: out_word = 8'h05;
		16'h33AD: out_word = 8'h00;
		16'h33AE: out_word = 8'hCD;
		16'h33AF: out_word = 8'h05;
		16'h33B0: out_word = 8'h1F;
		16'h33B1: out_word = 8'hE1;
		16'h33B2: out_word = 8'hD1;
		16'h33B3: out_word = 8'hC9;
		16'h33B4: out_word = 8'hED;
		16'h33B5: out_word = 8'h5B;
		16'h33B6: out_word = 8'h65;
		16'h33B7: out_word = 8'h5C;
		16'h33B8: out_word = 8'hCD;
		16'h33B9: out_word = 8'hC0;
		16'h33BA: out_word = 8'h33;
		16'h33BB: out_word = 8'hED;
		16'h33BC: out_word = 8'h53;
		16'h33BD: out_word = 8'h65;
		16'h33BE: out_word = 8'h5C;
		16'h33BF: out_word = 8'hC9;
		16'h33C0: out_word = 8'hCD;
		16'h33C1: out_word = 8'hA9;
		16'h33C2: out_word = 8'h33;
		16'h33C3: out_word = 8'hED;
		16'h33C4: out_word = 8'hB0;
		16'h33C5: out_word = 8'hC9;
		16'h33C6: out_word = 8'h62;
		16'h33C7: out_word = 8'h6B;
		16'h33C8: out_word = 8'hCD;
		16'h33C9: out_word = 8'hA9;
		16'h33CA: out_word = 8'h33;
		16'h33CB: out_word = 8'hD9;
		16'h33CC: out_word = 8'hE5;
		16'h33CD: out_word = 8'hD9;
		16'h33CE: out_word = 8'hE3;
		16'h33CF: out_word = 8'hC5;
		16'h33D0: out_word = 8'h7E;
		16'h33D1: out_word = 8'hE6;
		16'h33D2: out_word = 8'hC0;
		16'h33D3: out_word = 8'h07;
		16'h33D4: out_word = 8'h07;
		16'h33D5: out_word = 8'h4F;
		16'h33D6: out_word = 8'h0C;
		16'h33D7: out_word = 8'h7E;
		16'h33D8: out_word = 8'hE6;
		16'h33D9: out_word = 8'h3F;
		16'h33DA: out_word = 8'h20;
		16'h33DB: out_word = 8'h02;
		16'h33DC: out_word = 8'h23;
		16'h33DD: out_word = 8'h7E;
		16'h33DE: out_word = 8'hC6;
		16'h33DF: out_word = 8'h50;
		16'h33E0: out_word = 8'h12;
		16'h33E1: out_word = 8'h3E;
		16'h33E2: out_word = 8'h05;
		16'h33E3: out_word = 8'h91;
		16'h33E4: out_word = 8'h23;
		16'h33E5: out_word = 8'h13;
		16'h33E6: out_word = 8'h06;
		16'h33E7: out_word = 8'h00;
		16'h33E8: out_word = 8'hED;
		16'h33E9: out_word = 8'hB0;
		16'h33EA: out_word = 8'hC1;
		16'h33EB: out_word = 8'hE3;
		16'h33EC: out_word = 8'hD9;
		16'h33ED: out_word = 8'hE1;
		16'h33EE: out_word = 8'hD9;
		16'h33EF: out_word = 8'h47;
		16'h33F0: out_word = 8'hAF;
		16'h33F1: out_word = 8'h05;
		16'h33F2: out_word = 8'hC8;
		16'h33F3: out_word = 8'h12;
		16'h33F4: out_word = 8'h13;
		16'h33F5: out_word = 8'h18;
		16'h33F6: out_word = 8'hFA;
		16'h33F7: out_word = 8'hA7;
		16'h33F8: out_word = 8'hC8;
		16'h33F9: out_word = 8'hF5;
		16'h33FA: out_word = 8'hD5;
		16'h33FB: out_word = 8'h11;
		16'h33FC: out_word = 8'h00;
		16'h33FD: out_word = 8'h00;
		16'h33FE: out_word = 8'hCD;
		16'h33FF: out_word = 8'hC8;
		16'h3400: out_word = 8'h33;
		16'h3401: out_word = 8'hD1;
		16'h3402: out_word = 8'hF1;
		16'h3403: out_word = 8'h3D;
		16'h3404: out_word = 8'h18;
		16'h3405: out_word = 8'hF2;
		16'h3406: out_word = 8'h4F;
		16'h3407: out_word = 8'h07;
		16'h3408: out_word = 8'h07;
		16'h3409: out_word = 8'h81;
		16'h340A: out_word = 8'h4F;
		16'h340B: out_word = 8'h06;
		16'h340C: out_word = 8'h00;
		16'h340D: out_word = 8'h09;
		16'h340E: out_word = 8'hC9;
		16'h340F: out_word = 8'hD5;
		16'h3410: out_word = 8'h2A;
		16'h3411: out_word = 8'h68;
		16'h3412: out_word = 8'h5C;
		16'h3413: out_word = 8'hCD;
		16'h3414: out_word = 8'h06;
		16'h3415: out_word = 8'h34;
		16'h3416: out_word = 8'hCD;
		16'h3417: out_word = 8'hC0;
		16'h3418: out_word = 8'h33;
		16'h3419: out_word = 8'hE1;
		16'h341A: out_word = 8'hC9;
		16'h341B: out_word = 8'h62;
		16'h341C: out_word = 8'h6B;
		16'h341D: out_word = 8'hD9;
		16'h341E: out_word = 8'hE5;
		16'h341F: out_word = 8'h21;
		16'h3420: out_word = 8'hC5;
		16'h3421: out_word = 8'h32;
		16'h3422: out_word = 8'hD9;
		16'h3423: out_word = 8'hCD;
		16'h3424: out_word = 8'hF7;
		16'h3425: out_word = 8'h33;
		16'h3426: out_word = 8'hCD;
		16'h3427: out_word = 8'hC8;
		16'h3428: out_word = 8'h33;
		16'h3429: out_word = 8'hD9;
		16'h342A: out_word = 8'hE1;
		16'h342B: out_word = 8'hD9;
		16'h342C: out_word = 8'hC9;
		16'h342D: out_word = 8'hE5;
		16'h342E: out_word = 8'hEB;
		16'h342F: out_word = 8'h2A;
		16'h3430: out_word = 8'h68;
		16'h3431: out_word = 8'h5C;
		16'h3432: out_word = 8'hCD;
		16'h3433: out_word = 8'h06;
		16'h3434: out_word = 8'h34;
		16'h3435: out_word = 8'hEB;
		16'h3436: out_word = 8'hCD;
		16'h3437: out_word = 8'hC0;
		16'h3438: out_word = 8'h33;
		16'h3439: out_word = 8'hEB;
		16'h343A: out_word = 8'hE1;
		16'h343B: out_word = 8'hC9;
		16'h343C: out_word = 8'h06;
		16'h343D: out_word = 8'h05;
		16'h343E: out_word = 8'h1A;
		16'h343F: out_word = 8'h4E;
		16'h3440: out_word = 8'hEB;
		16'h3441: out_word = 8'h12;
		16'h3442: out_word = 8'h71;
		16'h3443: out_word = 8'h23;
		16'h3444: out_word = 8'h13;
		16'h3445: out_word = 8'h10;
		16'h3446: out_word = 8'hF7;
		16'h3447: out_word = 8'hEB;
		16'h3448: out_word = 8'hC9;
		16'h3449: out_word = 8'h47;
		16'h344A: out_word = 8'hCD;
		16'h344B: out_word = 8'h5E;
		16'h344C: out_word = 8'h33;
		16'h344D: out_word = 8'h31;
		16'h344E: out_word = 8'h0F;
		16'h344F: out_word = 8'hC0;
		16'h3450: out_word = 8'h02;
		16'h3451: out_word = 8'hA0;
		16'h3452: out_word = 8'hC2;
		16'h3453: out_word = 8'h31;
		16'h3454: out_word = 8'hE0;
		16'h3455: out_word = 8'h04;
		16'h3456: out_word = 8'hE2;
		16'h3457: out_word = 8'hC1;
		16'h3458: out_word = 8'h03;
		16'h3459: out_word = 8'h38;
		16'h345A: out_word = 8'hCD;
		16'h345B: out_word = 8'hC6;
		16'h345C: out_word = 8'h33;
		16'h345D: out_word = 8'hCD;
		16'h345E: out_word = 8'h62;
		16'h345F: out_word = 8'h33;
		16'h3460: out_word = 8'h0F;
		16'h3461: out_word = 8'h01;
		16'h3462: out_word = 8'hC2;
		16'h3463: out_word = 8'h02;
		16'h3464: out_word = 8'h35;
		16'h3465: out_word = 8'hEE;
		16'h3466: out_word = 8'hE1;
		16'h3467: out_word = 8'h03;
		16'h3468: out_word = 8'h38;
		16'h3469: out_word = 8'hC9;
		16'h346A: out_word = 8'h06;
		16'h346B: out_word = 8'hFF;
		16'h346C: out_word = 8'h18;
		16'h346D: out_word = 8'h06;
		16'h346E: out_word = 8'hCD;
		16'h346F: out_word = 8'hE9;
		16'h3470: out_word = 8'h34;
		16'h3471: out_word = 8'hD8;
		16'h3472: out_word = 8'h06;
		16'h3473: out_word = 8'h00;
		16'h3474: out_word = 8'h7E;
		16'h3475: out_word = 8'hA7;
		16'h3476: out_word = 8'h28;
		16'h3477: out_word = 8'h0B;
		16'h3478: out_word = 8'h23;
		16'h3479: out_word = 8'h78;
		16'h347A: out_word = 8'hE6;
		16'h347B: out_word = 8'h80;
		16'h347C: out_word = 8'hB6;
		16'h347D: out_word = 8'h17;
		16'h347E: out_word = 8'h3F;
		16'h347F: out_word = 8'h1F;
		16'h3480: out_word = 8'h77;
		16'h3481: out_word = 8'h2B;
		16'h3482: out_word = 8'hC9;
		16'h3483: out_word = 8'hD5;
		16'h3484: out_word = 8'hE5;
		16'h3485: out_word = 8'hCD;
		16'h3486: out_word = 8'h7F;
		16'h3487: out_word = 8'h2D;
		16'h3488: out_word = 8'hE1;
		16'h3489: out_word = 8'h78;
		16'h348A: out_word = 8'hB1;
		16'h348B: out_word = 8'h2F;
		16'h348C: out_word = 8'h4F;
		16'h348D: out_word = 8'hCD;
		16'h348E: out_word = 8'h8E;
		16'h348F: out_word = 8'h2D;
		16'h3490: out_word = 8'hD1;
		16'h3491: out_word = 8'hC9;
		16'h3492: out_word = 8'hCD;
		16'h3493: out_word = 8'hE9;
		16'h3494: out_word = 8'h34;
		16'h3495: out_word = 8'hD8;
		16'h3496: out_word = 8'hD5;
		16'h3497: out_word = 8'h11;
		16'h3498: out_word = 8'h01;
		16'h3499: out_word = 8'h00;
		16'h349A: out_word = 8'h23;
		16'h349B: out_word = 8'hCB;
		16'h349C: out_word = 8'h16;
		16'h349D: out_word = 8'h2B;
		16'h349E: out_word = 8'h9F;
		16'h349F: out_word = 8'h4F;
		16'h34A0: out_word = 8'hCD;
		16'h34A1: out_word = 8'h8E;
		16'h34A2: out_word = 8'h2D;
		16'h34A3: out_word = 8'hD1;
		16'h34A4: out_word = 8'hC9;
		16'h34A5: out_word = 8'hCD;
		16'h34A6: out_word = 8'h99;
		16'h34A7: out_word = 8'h1E;
		16'h34A8: out_word = 8'hED;
		16'h34A9: out_word = 8'h78;
		16'h34AA: out_word = 8'h18;
		16'h34AB: out_word = 8'h04;
		16'h34AC: out_word = 8'hCD;
		16'h34AD: out_word = 8'h99;
		16'h34AE: out_word = 8'h1E;
		16'h34AF: out_word = 8'h0A;
		16'h34B0: out_word = 8'hC3;
		16'h34B1: out_word = 8'h28;
		16'h34B2: out_word = 8'h2D;
		16'h34B3: out_word = 8'hCD;
		16'h34B4: out_word = 8'h99;
		16'h34B5: out_word = 8'h1E;
		16'h34B6: out_word = 8'h21;
		16'h34B7: out_word = 8'h2B;
		16'h34B8: out_word = 8'h2D;
		16'h34B9: out_word = 8'hE5;
		16'h34BA: out_word = 8'hC5;
		16'h34BB: out_word = 8'hC9;
		16'h34BC: out_word = 8'hCD;
		16'h34BD: out_word = 8'hF1;
		16'h34BE: out_word = 8'h2B;
		16'h34BF: out_word = 8'h0B;
		16'h34C0: out_word = 8'h78;
		16'h34C1: out_word = 8'hB1;
		16'h34C2: out_word = 8'h20;
		16'h34C3: out_word = 8'h23;
		16'h34C4: out_word = 8'h1A;
		16'h34C5: out_word = 8'hCD;
		16'h34C6: out_word = 8'h8D;
		16'h34C7: out_word = 8'h2C;
		16'h34C8: out_word = 8'h38;
		16'h34C9: out_word = 8'h09;
		16'h34CA: out_word = 8'hD6;
		16'h34CB: out_word = 8'h90;
		16'h34CC: out_word = 8'h38;
		16'h34CD: out_word = 8'h19;
		16'h34CE: out_word = 8'hFE;
		16'h34CF: out_word = 8'h15;
		16'h34D0: out_word = 8'h30;
		16'h34D1: out_word = 8'h15;
		16'h34D2: out_word = 8'h3C;
		16'h34D3: out_word = 8'h3D;
		16'h34D4: out_word = 8'h87;
		16'h34D5: out_word = 8'h87;
		16'h34D6: out_word = 8'h87;
		16'h34D7: out_word = 8'hFE;
		16'h34D8: out_word = 8'hA8;
		16'h34D9: out_word = 8'h30;
		16'h34DA: out_word = 8'h0C;
		16'h34DB: out_word = 8'hED;
		16'h34DC: out_word = 8'h4B;
		16'h34DD: out_word = 8'h7B;
		16'h34DE: out_word = 8'h5C;
		16'h34DF: out_word = 8'h81;
		16'h34E0: out_word = 8'h4F;
		16'h34E1: out_word = 8'h30;
		16'h34E2: out_word = 8'h01;
		16'h34E3: out_word = 8'h04;
		16'h34E4: out_word = 8'hC3;
		16'h34E5: out_word = 8'h2B;
		16'h34E6: out_word = 8'h2D;
		16'h34E7: out_word = 8'hCF;
		16'h34E8: out_word = 8'h09;
		16'h34E9: out_word = 8'hE5;
		16'h34EA: out_word = 8'hC5;
		16'h34EB: out_word = 8'h47;
		16'h34EC: out_word = 8'h7E;
		16'h34ED: out_word = 8'h23;
		16'h34EE: out_word = 8'hB6;
		16'h34EF: out_word = 8'h23;
		16'h34F0: out_word = 8'hB6;
		16'h34F1: out_word = 8'h23;
		16'h34F2: out_word = 8'hB6;
		16'h34F3: out_word = 8'h78;
		16'h34F4: out_word = 8'hC1;
		16'h34F5: out_word = 8'hE1;
		16'h34F6: out_word = 8'hC0;
		16'h34F7: out_word = 8'h37;
		16'h34F8: out_word = 8'hC9;
		16'h34F9: out_word = 8'hCD;
		16'h34FA: out_word = 8'hE9;
		16'h34FB: out_word = 8'h34;
		16'h34FC: out_word = 8'hD8;
		16'h34FD: out_word = 8'h3E;
		16'h34FE: out_word = 8'hFF;
		16'h34FF: out_word = 8'h18;
		16'h3500: out_word = 8'h06;
		16'h3501: out_word = 8'hCD;
		16'h3502: out_word = 8'hE9;
		16'h3503: out_word = 8'h34;
		16'h3504: out_word = 8'h18;
		16'h3505: out_word = 8'h05;
		16'h3506: out_word = 8'hAF;
		16'h3507: out_word = 8'h23;
		16'h3508: out_word = 8'hAE;
		16'h3509: out_word = 8'h2B;
		16'h350A: out_word = 8'h07;
		16'h350B: out_word = 8'hE5;
		16'h350C: out_word = 8'h3E;
		16'h350D: out_word = 8'h00;
		16'h350E: out_word = 8'h77;
		16'h350F: out_word = 8'h23;
		16'h3510: out_word = 8'h77;
		16'h3511: out_word = 8'h23;
		16'h3512: out_word = 8'h17;
		16'h3513: out_word = 8'h77;
		16'h3514: out_word = 8'h1F;
		16'h3515: out_word = 8'h23;
		16'h3516: out_word = 8'h77;
		16'h3517: out_word = 8'h23;
		16'h3518: out_word = 8'h77;
		16'h3519: out_word = 8'hE1;
		16'h351A: out_word = 8'hC9;
		16'h351B: out_word = 8'hEB;
		16'h351C: out_word = 8'hCD;
		16'h351D: out_word = 8'hE9;
		16'h351E: out_word = 8'h34;
		16'h351F: out_word = 8'hEB;
		16'h3520: out_word = 8'hD8;
		16'h3521: out_word = 8'h37;
		16'h3522: out_word = 8'h18;
		16'h3523: out_word = 8'hE7;
		16'h3524: out_word = 8'hEB;
		16'h3525: out_word = 8'hCD;
		16'h3526: out_word = 8'hE9;
		16'h3527: out_word = 8'h34;
		16'h3528: out_word = 8'hEB;
		16'h3529: out_word = 8'hD0;
		16'h352A: out_word = 8'hA7;
		16'h352B: out_word = 8'h18;
		16'h352C: out_word = 8'hDE;
		16'h352D: out_word = 8'hEB;
		16'h352E: out_word = 8'hCD;
		16'h352F: out_word = 8'hE9;
		16'h3530: out_word = 8'h34;
		16'h3531: out_word = 8'hEB;
		16'h3532: out_word = 8'hD0;
		16'h3533: out_word = 8'hD5;
		16'h3534: out_word = 8'h1B;
		16'h3535: out_word = 8'hAF;
		16'h3536: out_word = 8'h12;
		16'h3537: out_word = 8'h1B;
		16'h3538: out_word = 8'h12;
		16'h3539: out_word = 8'hD1;
		16'h353A: out_word = 8'hC9;
		16'h353B: out_word = 8'h78;
		16'h353C: out_word = 8'hD6;
		16'h353D: out_word = 8'h08;
		16'h353E: out_word = 8'hCB;
		16'h353F: out_word = 8'h57;
		16'h3540: out_word = 8'h20;
		16'h3541: out_word = 8'h01;
		16'h3542: out_word = 8'h3D;
		16'h3543: out_word = 8'h0F;
		16'h3544: out_word = 8'h30;
		16'h3545: out_word = 8'h08;
		16'h3546: out_word = 8'hF5;
		16'h3547: out_word = 8'hE5;
		16'h3548: out_word = 8'hCD;
		16'h3549: out_word = 8'h3C;
		16'h354A: out_word = 8'h34;
		16'h354B: out_word = 8'hD1;
		16'h354C: out_word = 8'hEB;
		16'h354D: out_word = 8'hF1;
		16'h354E: out_word = 8'hCB;
		16'h354F: out_word = 8'h57;
		16'h3550: out_word = 8'h20;
		16'h3551: out_word = 8'h07;
		16'h3552: out_word = 8'h0F;
		16'h3553: out_word = 8'hF5;
		16'h3554: out_word = 8'hCD;
		16'h3555: out_word = 8'h0F;
		16'h3556: out_word = 8'h30;
		16'h3557: out_word = 8'h18;
		16'h3558: out_word = 8'h33;
		16'h3559: out_word = 8'h0F;
		16'h355A: out_word = 8'hF5;
		16'h355B: out_word = 8'hCD;
		16'h355C: out_word = 8'hF1;
		16'h355D: out_word = 8'h2B;
		16'h355E: out_word = 8'hD5;
		16'h355F: out_word = 8'hC5;
		16'h3560: out_word = 8'hCD;
		16'h3561: out_word = 8'hF1;
		16'h3562: out_word = 8'h2B;
		16'h3563: out_word = 8'hE1;
		16'h3564: out_word = 8'h7C;
		16'h3565: out_word = 8'hB5;
		16'h3566: out_word = 8'hE3;
		16'h3567: out_word = 8'h78;
		16'h3568: out_word = 8'h20;
		16'h3569: out_word = 8'h0B;
		16'h356A: out_word = 8'hB1;
		16'h356B: out_word = 8'hC1;
		16'h356C: out_word = 8'h28;
		16'h356D: out_word = 8'h04;
		16'h356E: out_word = 8'hF1;
		16'h356F: out_word = 8'h3F;
		16'h3570: out_word = 8'h18;
		16'h3571: out_word = 8'h16;
		16'h3572: out_word = 8'hF1;
		16'h3573: out_word = 8'h18;
		16'h3574: out_word = 8'h13;
		16'h3575: out_word = 8'hB1;
		16'h3576: out_word = 8'h28;
		16'h3577: out_word = 8'h0D;
		16'h3578: out_word = 8'h1A;
		16'h3579: out_word = 8'h96;
		16'h357A: out_word = 8'h38;
		16'h357B: out_word = 8'h09;
		16'h357C: out_word = 8'h20;
		16'h357D: out_word = 8'hED;
		16'h357E: out_word = 8'h0B;
		16'h357F: out_word = 8'h13;
		16'h3580: out_word = 8'h23;
		16'h3581: out_word = 8'hE3;
		16'h3582: out_word = 8'h2B;
		16'h3583: out_word = 8'h18;
		16'h3584: out_word = 8'hDF;
		16'h3585: out_word = 8'hC1;
		16'h3586: out_word = 8'hF1;
		16'h3587: out_word = 8'hA7;
		16'h3588: out_word = 8'hF5;
		16'h3589: out_word = 8'hEF;
		16'h358A: out_word = 8'hA0;
		16'h358B: out_word = 8'h38;
		16'h358C: out_word = 8'hF1;
		16'h358D: out_word = 8'hF5;
		16'h358E: out_word = 8'hDC;
		16'h358F: out_word = 8'h01;
		16'h3590: out_word = 8'h35;
		16'h3591: out_word = 8'hF1;
		16'h3592: out_word = 8'hF5;
		16'h3593: out_word = 8'hD4;
		16'h3594: out_word = 8'hF9;
		16'h3595: out_word = 8'h34;
		16'h3596: out_word = 8'hF1;
		16'h3597: out_word = 8'h0F;
		16'h3598: out_word = 8'hD4;
		16'h3599: out_word = 8'h01;
		16'h359A: out_word = 8'h35;
		16'h359B: out_word = 8'hC9;
		16'h359C: out_word = 8'hCD;
		16'h359D: out_word = 8'hF1;
		16'h359E: out_word = 8'h2B;
		16'h359F: out_word = 8'hD5;
		16'h35A0: out_word = 8'hC5;
		16'h35A1: out_word = 8'hCD;
		16'h35A2: out_word = 8'hF1;
		16'h35A3: out_word = 8'h2B;
		16'h35A4: out_word = 8'hE1;
		16'h35A5: out_word = 8'hE5;
		16'h35A6: out_word = 8'hD5;
		16'h35A7: out_word = 8'hC5;
		16'h35A8: out_word = 8'h09;
		16'h35A9: out_word = 8'h44;
		16'h35AA: out_word = 8'h4D;
		16'h35AB: out_word = 8'hF7;
		16'h35AC: out_word = 8'hCD;
		16'h35AD: out_word = 8'hB2;
		16'h35AE: out_word = 8'h2A;
		16'h35AF: out_word = 8'hC1;
		16'h35B0: out_word = 8'hE1;
		16'h35B1: out_word = 8'h78;
		16'h35B2: out_word = 8'hB1;
		16'h35B3: out_word = 8'h28;
		16'h35B4: out_word = 8'h02;
		16'h35B5: out_word = 8'hED;
		16'h35B6: out_word = 8'hB0;
		16'h35B7: out_word = 8'hC1;
		16'h35B8: out_word = 8'hE1;
		16'h35B9: out_word = 8'h78;
		16'h35BA: out_word = 8'hB1;
		16'h35BB: out_word = 8'h28;
		16'h35BC: out_word = 8'h02;
		16'h35BD: out_word = 8'hED;
		16'h35BE: out_word = 8'hB0;
		16'h35BF: out_word = 8'h2A;
		16'h35C0: out_word = 8'h65;
		16'h35C1: out_word = 8'h5C;
		16'h35C2: out_word = 8'h11;
		16'h35C3: out_word = 8'hFB;
		16'h35C4: out_word = 8'hFF;
		16'h35C5: out_word = 8'hE5;
		16'h35C6: out_word = 8'h19;
		16'h35C7: out_word = 8'hD1;
		16'h35C8: out_word = 8'hC9;
		16'h35C9: out_word = 8'hCD;
		16'h35CA: out_word = 8'hD5;
		16'h35CB: out_word = 8'h2D;
		16'h35CC: out_word = 8'h38;
		16'h35CD: out_word = 8'h0E;
		16'h35CE: out_word = 8'h20;
		16'h35CF: out_word = 8'h0C;
		16'h35D0: out_word = 8'hF5;
		16'h35D1: out_word = 8'h01;
		16'h35D2: out_word = 8'h01;
		16'h35D3: out_word = 8'h00;
		16'h35D4: out_word = 8'hF7;
		16'h35D5: out_word = 8'hF1;
		16'h35D6: out_word = 8'h12;
		16'h35D7: out_word = 8'hCD;
		16'h35D8: out_word = 8'hB2;
		16'h35D9: out_word = 8'h2A;
		16'h35DA: out_word = 8'hEB;
		16'h35DB: out_word = 8'hC9;
		16'h35DC: out_word = 8'hCF;
		16'h35DD: out_word = 8'h0A;
		16'h35DE: out_word = 8'h2A;
		16'h35DF: out_word = 8'h5D;
		16'h35E0: out_word = 8'h5C;
		16'h35E1: out_word = 8'hE5;
		16'h35E2: out_word = 8'h78;
		16'h35E3: out_word = 8'hC6;
		16'h35E4: out_word = 8'hE3;
		16'h35E5: out_word = 8'h9F;
		16'h35E6: out_word = 8'hF5;
		16'h35E7: out_word = 8'hCD;
		16'h35E8: out_word = 8'hF1;
		16'h35E9: out_word = 8'h2B;
		16'h35EA: out_word = 8'hD5;
		16'h35EB: out_word = 8'h03;
		16'h35EC: out_word = 8'hF7;
		16'h35ED: out_word = 8'hE1;
		16'h35EE: out_word = 8'hED;
		16'h35EF: out_word = 8'h53;
		16'h35F0: out_word = 8'h5D;
		16'h35F1: out_word = 8'h5C;
		16'h35F2: out_word = 8'hD5;
		16'h35F3: out_word = 8'hED;
		16'h35F4: out_word = 8'hB0;
		16'h35F5: out_word = 8'hEB;
		16'h35F6: out_word = 8'h2B;
		16'h35F7: out_word = 8'h36;
		16'h35F8: out_word = 8'h0D;
		16'h35F9: out_word = 8'hFD;
		16'h35FA: out_word = 8'hCB;
		16'h35FB: out_word = 8'h01;
		16'h35FC: out_word = 8'hBE;
		16'h35FD: out_word = 8'hCD;
		16'h35FE: out_word = 8'hFB;
		16'h35FF: out_word = 8'h24;
		16'h3600: out_word = 8'hDF;
		16'h3601: out_word = 8'hFE;
		16'h3602: out_word = 8'h0D;
		16'h3603: out_word = 8'h20;
		16'h3604: out_word = 8'h07;
		16'h3605: out_word = 8'hE1;
		16'h3606: out_word = 8'hF1;
		16'h3607: out_word = 8'hFD;
		16'h3608: out_word = 8'hAE;
		16'h3609: out_word = 8'h01;
		16'h360A: out_word = 8'hE6;
		16'h360B: out_word = 8'h40;
		16'h360C: out_word = 8'hC2;
		16'h360D: out_word = 8'h8A;
		16'h360E: out_word = 8'h1C;
		16'h360F: out_word = 8'h22;
		16'h3610: out_word = 8'h5D;
		16'h3611: out_word = 8'h5C;
		16'h3612: out_word = 8'hFD;
		16'h3613: out_word = 8'hCB;
		16'h3614: out_word = 8'h01;
		16'h3615: out_word = 8'hFE;
		16'h3616: out_word = 8'hCD;
		16'h3617: out_word = 8'hFB;
		16'h3618: out_word = 8'h24;
		16'h3619: out_word = 8'hE1;
		16'h361A: out_word = 8'h22;
		16'h361B: out_word = 8'h5D;
		16'h361C: out_word = 8'h5C;
		16'h361D: out_word = 8'h18;
		16'h361E: out_word = 8'hA0;
		16'h361F: out_word = 8'h01;
		16'h3620: out_word = 8'h01;
		16'h3621: out_word = 8'h00;
		16'h3622: out_word = 8'hF7;
		16'h3623: out_word = 8'h22;
		16'h3624: out_word = 8'h5B;
		16'h3625: out_word = 8'h5C;
		16'h3626: out_word = 8'hE5;
		16'h3627: out_word = 8'h2A;
		16'h3628: out_word = 8'h51;
		16'h3629: out_word = 8'h5C;
		16'h362A: out_word = 8'hE5;
		16'h362B: out_word = 8'h3E;
		16'h362C: out_word = 8'hFF;
		16'h362D: out_word = 8'hCD;
		16'h362E: out_word = 8'h01;
		16'h362F: out_word = 8'h16;
		16'h3630: out_word = 8'hCD;
		16'h3631: out_word = 8'hE3;
		16'h3632: out_word = 8'h2D;
		16'h3633: out_word = 8'hE1;
		16'h3634: out_word = 8'hCD;
		16'h3635: out_word = 8'h15;
		16'h3636: out_word = 8'h16;
		16'h3637: out_word = 8'hD1;
		16'h3638: out_word = 8'h2A;
		16'h3639: out_word = 8'h5B;
		16'h363A: out_word = 8'h5C;
		16'h363B: out_word = 8'hA7;
		16'h363C: out_word = 8'hED;
		16'h363D: out_word = 8'h52;
		16'h363E: out_word = 8'h44;
		16'h363F: out_word = 8'h4D;
		16'h3640: out_word = 8'hCD;
		16'h3641: out_word = 8'hB2;
		16'h3642: out_word = 8'h2A;
		16'h3643: out_word = 8'hEB;
		16'h3644: out_word = 8'hC9;
		16'h3645: out_word = 8'hCD;
		16'h3646: out_word = 8'h94;
		16'h3647: out_word = 8'h1E;
		16'h3648: out_word = 8'hFE;
		16'h3649: out_word = 8'h10;
		16'h364A: out_word = 8'hD2;
		16'h364B: out_word = 8'h9F;
		16'h364C: out_word = 8'h1E;
		16'h364D: out_word = 8'h2A;
		16'h364E: out_word = 8'h51;
		16'h364F: out_word = 8'h5C;
		16'h3650: out_word = 8'hE5;
		16'h3651: out_word = 8'hCD;
		16'h3652: out_word = 8'h01;
		16'h3653: out_word = 8'h16;
		16'h3654: out_word = 8'hCD;
		16'h3655: out_word = 8'hE6;
		16'h3656: out_word = 8'h15;
		16'h3657: out_word = 8'h01;
		16'h3658: out_word = 8'h00;
		16'h3659: out_word = 8'h00;
		16'h365A: out_word = 8'h30;
		16'h365B: out_word = 8'h03;
		16'h365C: out_word = 8'h0C;
		16'h365D: out_word = 8'hF7;
		16'h365E: out_word = 8'h12;
		16'h365F: out_word = 8'hCD;
		16'h3660: out_word = 8'hB2;
		16'h3661: out_word = 8'h2A;
		16'h3662: out_word = 8'hE1;
		16'h3663: out_word = 8'hCD;
		16'h3664: out_word = 8'h15;
		16'h3665: out_word = 8'h16;
		16'h3666: out_word = 8'hC3;
		16'h3667: out_word = 8'hBF;
		16'h3668: out_word = 8'h35;
		16'h3669: out_word = 8'hCD;
		16'h366A: out_word = 8'hF1;
		16'h366B: out_word = 8'h2B;
		16'h366C: out_word = 8'h78;
		16'h366D: out_word = 8'hB1;
		16'h366E: out_word = 8'h28;
		16'h366F: out_word = 8'h01;
		16'h3670: out_word = 8'h1A;
		16'h3671: out_word = 8'hC3;
		16'h3672: out_word = 8'h28;
		16'h3673: out_word = 8'h2D;
		16'h3674: out_word = 8'hCD;
		16'h3675: out_word = 8'hF1;
		16'h3676: out_word = 8'h2B;
		16'h3677: out_word = 8'hC3;
		16'h3678: out_word = 8'h2B;
		16'h3679: out_word = 8'h2D;
		16'h367A: out_word = 8'hD9;
		16'h367B: out_word = 8'hE5;
		16'h367C: out_word = 8'h21;
		16'h367D: out_word = 8'h67;
		16'h367E: out_word = 8'h5C;
		16'h367F: out_word = 8'h35;
		16'h3680: out_word = 8'hE1;
		16'h3681: out_word = 8'h20;
		16'h3682: out_word = 8'h04;
		16'h3683: out_word = 8'h23;
		16'h3684: out_word = 8'hD9;
		16'h3685: out_word = 8'hC9;
		16'h3686: out_word = 8'hD9;
		16'h3687: out_word = 8'h5E;
		16'h3688: out_word = 8'h7B;
		16'h3689: out_word = 8'h17;
		16'h368A: out_word = 8'h9F;
		16'h368B: out_word = 8'h57;
		16'h368C: out_word = 8'h19;
		16'h368D: out_word = 8'hD9;
		16'h368E: out_word = 8'hC9;
		16'h368F: out_word = 8'h13;
		16'h3690: out_word = 8'h13;
		16'h3691: out_word = 8'h1A;
		16'h3692: out_word = 8'h1B;
		16'h3693: out_word = 8'h1B;
		16'h3694: out_word = 8'hA7;
		16'h3695: out_word = 8'h20;
		16'h3696: out_word = 8'hEF;
		16'h3697: out_word = 8'hD9;
		16'h3698: out_word = 8'h23;
		16'h3699: out_word = 8'hD9;
		16'h369A: out_word = 8'hC9;
		16'h369B: out_word = 8'hF1;
		16'h369C: out_word = 8'hD9;
		16'h369D: out_word = 8'hE3;
		16'h369E: out_word = 8'hD9;
		16'h369F: out_word = 8'hC9;
		16'h36A0: out_word = 8'hEF;
		16'h36A1: out_word = 8'hC0;
		16'h36A2: out_word = 8'h02;
		16'h36A3: out_word = 8'h31;
		16'h36A4: out_word = 8'hE0;
		16'h36A5: out_word = 8'h05;
		16'h36A6: out_word = 8'h27;
		16'h36A7: out_word = 8'hE0;
		16'h36A8: out_word = 8'h01;
		16'h36A9: out_word = 8'hC0;
		16'h36AA: out_word = 8'h04;
		16'h36AB: out_word = 8'h03;
		16'h36AC: out_word = 8'hE0;
		16'h36AD: out_word = 8'h38;
		16'h36AE: out_word = 8'hC9;
		16'h36AF: out_word = 8'hEF;
		16'h36B0: out_word = 8'h31;
		16'h36B1: out_word = 8'h36;
		16'h36B2: out_word = 8'h00;
		16'h36B3: out_word = 8'h04;
		16'h36B4: out_word = 8'h3A;
		16'h36B5: out_word = 8'h38;
		16'h36B6: out_word = 8'hC9;
		16'h36B7: out_word = 8'h31;
		16'h36B8: out_word = 8'h3A;
		16'h36B9: out_word = 8'hC0;
		16'h36BA: out_word = 8'h03;
		16'h36BB: out_word = 8'hE0;
		16'h36BC: out_word = 8'h01;
		16'h36BD: out_word = 8'h30;
		16'h36BE: out_word = 8'h00;
		16'h36BF: out_word = 8'h03;
		16'h36C0: out_word = 8'hA1;
		16'h36C1: out_word = 8'h03;
		16'h36C2: out_word = 8'h38;
		16'h36C3: out_word = 8'hC9;
		16'h36C4: out_word = 8'hEF;
		16'h36C5: out_word = 8'h3D;
		16'h36C6: out_word = 8'h34;
		16'h36C7: out_word = 8'hF1;
		16'h36C8: out_word = 8'h38;
		16'h36C9: out_word = 8'hAA;
		16'h36CA: out_word = 8'h3B;
		16'h36CB: out_word = 8'h29;
		16'h36CC: out_word = 8'h04;
		16'h36CD: out_word = 8'h31;
		16'h36CE: out_word = 8'h27;
		16'h36CF: out_word = 8'hC3;
		16'h36D0: out_word = 8'h03;
		16'h36D1: out_word = 8'h31;
		16'h36D2: out_word = 8'h0F;
		16'h36D3: out_word = 8'hA1;
		16'h36D4: out_word = 8'h03;
		16'h36D5: out_word = 8'h88;
		16'h36D6: out_word = 8'h13;
		16'h36D7: out_word = 8'h36;
		16'h36D8: out_word = 8'h58;
		16'h36D9: out_word = 8'h65;
		16'h36DA: out_word = 8'h66;
		16'h36DB: out_word = 8'h9D;
		16'h36DC: out_word = 8'h78;
		16'h36DD: out_word = 8'h65;
		16'h36DE: out_word = 8'h40;
		16'h36DF: out_word = 8'hA2;
		16'h36E0: out_word = 8'h60;
		16'h36E1: out_word = 8'h32;
		16'h36E2: out_word = 8'hC9;
		16'h36E3: out_word = 8'hE7;
		16'h36E4: out_word = 8'h21;
		16'h36E5: out_word = 8'hF7;
		16'h36E6: out_word = 8'hAF;
		16'h36E7: out_word = 8'h24;
		16'h36E8: out_word = 8'hEB;
		16'h36E9: out_word = 8'h2F;
		16'h36EA: out_word = 8'hB0;
		16'h36EB: out_word = 8'hB0;
		16'h36EC: out_word = 8'h14;
		16'h36ED: out_word = 8'hEE;
		16'h36EE: out_word = 8'h7E;
		16'h36EF: out_word = 8'hBB;
		16'h36F0: out_word = 8'h94;
		16'h36F1: out_word = 8'h58;
		16'h36F2: out_word = 8'hF1;
		16'h36F3: out_word = 8'h3A;
		16'h36F4: out_word = 8'h7E;
		16'h36F5: out_word = 8'hF8;
		16'h36F6: out_word = 8'hCF;
		16'h36F7: out_word = 8'hE3;
		16'h36F8: out_word = 8'h38;
		16'h36F9: out_word = 8'hCD;
		16'h36FA: out_word = 8'hD5;
		16'h36FB: out_word = 8'h2D;
		16'h36FC: out_word = 8'h20;
		16'h36FD: out_word = 8'h07;
		16'h36FE: out_word = 8'h38;
		16'h36FF: out_word = 8'h03;
		16'h3700: out_word = 8'h86;
		16'h3701: out_word = 8'h30;
		16'h3702: out_word = 8'h09;
		16'h3703: out_word = 8'hCF;
		16'h3704: out_word = 8'h05;
		16'h3705: out_word = 8'h38;
		16'h3706: out_word = 8'h07;
		16'h3707: out_word = 8'h96;
		16'h3708: out_word = 8'h30;
		16'h3709: out_word = 8'h04;
		16'h370A: out_word = 8'hED;
		16'h370B: out_word = 8'h44;
		16'h370C: out_word = 8'h77;
		16'h370D: out_word = 8'hC9;
		16'h370E: out_word = 8'hEF;
		16'h370F: out_word = 8'h02;
		16'h3710: out_word = 8'hA0;
		16'h3711: out_word = 8'h38;
		16'h3712: out_word = 8'hC9;
		16'h3713: out_word = 8'hEF;
		16'h3714: out_word = 8'h3D;
		16'h3715: out_word = 8'h31;
		16'h3716: out_word = 8'h37;
		16'h3717: out_word = 8'h00;
		16'h3718: out_word = 8'h04;
		16'h3719: out_word = 8'h38;
		16'h371A: out_word = 8'hCF;
		16'h371B: out_word = 8'h09;
		16'h371C: out_word = 8'hA0;
		16'h371D: out_word = 8'h02;
		16'h371E: out_word = 8'h38;
		16'h371F: out_word = 8'h7E;
		16'h3720: out_word = 8'h36;
		16'h3721: out_word = 8'h80;
		16'h3722: out_word = 8'hCD;
		16'h3723: out_word = 8'h28;
		16'h3724: out_word = 8'h2D;
		16'h3725: out_word = 8'hEF;
		16'h3726: out_word = 8'h34;
		16'h3727: out_word = 8'h38;
		16'h3728: out_word = 8'h00;
		16'h3729: out_word = 8'h03;
		16'h372A: out_word = 8'h01;
		16'h372B: out_word = 8'h31;
		16'h372C: out_word = 8'h34;
		16'h372D: out_word = 8'hF0;
		16'h372E: out_word = 8'h4C;
		16'h372F: out_word = 8'hCC;
		16'h3730: out_word = 8'hCC;
		16'h3731: out_word = 8'hCD;
		16'h3732: out_word = 8'h03;
		16'h3733: out_word = 8'h37;
		16'h3734: out_word = 8'h00;
		16'h3735: out_word = 8'h08;
		16'h3736: out_word = 8'h01;
		16'h3737: out_word = 8'hA1;
		16'h3738: out_word = 8'h03;
		16'h3739: out_word = 8'h01;
		16'h373A: out_word = 8'h38;
		16'h373B: out_word = 8'h34;
		16'h373C: out_word = 8'hEF;
		16'h373D: out_word = 8'h01;
		16'h373E: out_word = 8'h34;
		16'h373F: out_word = 8'hF0;
		16'h3740: out_word = 8'h31;
		16'h3741: out_word = 8'h72;
		16'h3742: out_word = 8'h17;
		16'h3743: out_word = 8'hF8;
		16'h3744: out_word = 8'h04;
		16'h3745: out_word = 8'h01;
		16'h3746: out_word = 8'hA2;
		16'h3747: out_word = 8'h03;
		16'h3748: out_word = 8'hA2;
		16'h3749: out_word = 8'h03;
		16'h374A: out_word = 8'h31;
		16'h374B: out_word = 8'h34;
		16'h374C: out_word = 8'h32;
		16'h374D: out_word = 8'h20;
		16'h374E: out_word = 8'h04;
		16'h374F: out_word = 8'hA2;
		16'h3750: out_word = 8'h03;
		16'h3751: out_word = 8'h8C;
		16'h3752: out_word = 8'h11;
		16'h3753: out_word = 8'hAC;
		16'h3754: out_word = 8'h14;
		16'h3755: out_word = 8'h09;
		16'h3756: out_word = 8'h56;
		16'h3757: out_word = 8'hDA;
		16'h3758: out_word = 8'hA5;
		16'h3759: out_word = 8'h59;
		16'h375A: out_word = 8'h30;
		16'h375B: out_word = 8'hC5;
		16'h375C: out_word = 8'h5C;
		16'h375D: out_word = 8'h90;
		16'h375E: out_word = 8'hAA;
		16'h375F: out_word = 8'h9E;
		16'h3760: out_word = 8'h70;
		16'h3761: out_word = 8'h6F;
		16'h3762: out_word = 8'h61;
		16'h3763: out_word = 8'hA1;
		16'h3764: out_word = 8'hCB;
		16'h3765: out_word = 8'hDA;
		16'h3766: out_word = 8'h96;
		16'h3767: out_word = 8'hA4;
		16'h3768: out_word = 8'h31;
		16'h3769: out_word = 8'h9F;
		16'h376A: out_word = 8'hB4;
		16'h376B: out_word = 8'hE7;
		16'h376C: out_word = 8'hA0;
		16'h376D: out_word = 8'hFE;
		16'h376E: out_word = 8'h5C;
		16'h376F: out_word = 8'hFC;
		16'h3770: out_word = 8'hEA;
		16'h3771: out_word = 8'h1B;
		16'h3772: out_word = 8'h43;
		16'h3773: out_word = 8'hCA;
		16'h3774: out_word = 8'h36;
		16'h3775: out_word = 8'hED;
		16'h3776: out_word = 8'hA7;
		16'h3777: out_word = 8'h9C;
		16'h3778: out_word = 8'h7E;
		16'h3779: out_word = 8'h5E;
		16'h377A: out_word = 8'hF0;
		16'h377B: out_word = 8'h6E;
		16'h377C: out_word = 8'h23;
		16'h377D: out_word = 8'h80;
		16'h377E: out_word = 8'h93;
		16'h377F: out_word = 8'h04;
		16'h3780: out_word = 8'h0F;
		16'h3781: out_word = 8'h38;
		16'h3782: out_word = 8'hC9;
		16'h3783: out_word = 8'hEF;
		16'h3784: out_word = 8'h3D;
		16'h3785: out_word = 8'h34;
		16'h3786: out_word = 8'hEE;
		16'h3787: out_word = 8'h22;
		16'h3788: out_word = 8'hF9;
		16'h3789: out_word = 8'h83;
		16'h378A: out_word = 8'h6E;
		16'h378B: out_word = 8'h04;
		16'h378C: out_word = 8'h31;
		16'h378D: out_word = 8'hA2;
		16'h378E: out_word = 8'h0F;
		16'h378F: out_word = 8'h27;
		16'h3790: out_word = 8'h03;
		16'h3791: out_word = 8'h31;
		16'h3792: out_word = 8'h0F;
		16'h3793: out_word = 8'h31;
		16'h3794: out_word = 8'h0F;
		16'h3795: out_word = 8'h31;
		16'h3796: out_word = 8'h2A;
		16'h3797: out_word = 8'hA1;
		16'h3798: out_word = 8'h03;
		16'h3799: out_word = 8'h31;
		16'h379A: out_word = 8'h37;
		16'h379B: out_word = 8'hC0;
		16'h379C: out_word = 8'h00;
		16'h379D: out_word = 8'h04;
		16'h379E: out_word = 8'h02;
		16'h379F: out_word = 8'h38;
		16'h37A0: out_word = 8'hC9;
		16'h37A1: out_word = 8'hA1;
		16'h37A2: out_word = 8'h03;
		16'h37A3: out_word = 8'h01;
		16'h37A4: out_word = 8'h36;
		16'h37A5: out_word = 8'h00;
		16'h37A6: out_word = 8'h02;
		16'h37A7: out_word = 8'h1B;
		16'h37A8: out_word = 8'h38;
		16'h37A9: out_word = 8'hC9;
		16'h37AA: out_word = 8'hEF;
		16'h37AB: out_word = 8'h39;
		16'h37AC: out_word = 8'h2A;
		16'h37AD: out_word = 8'hA1;
		16'h37AE: out_word = 8'h03;
		16'h37AF: out_word = 8'hE0;
		16'h37B0: out_word = 8'h00;
		16'h37B1: out_word = 8'h06;
		16'h37B2: out_word = 8'h1B;
		16'h37B3: out_word = 8'h33;
		16'h37B4: out_word = 8'h03;
		16'h37B5: out_word = 8'hEF;
		16'h37B6: out_word = 8'h39;
		16'h37B7: out_word = 8'h31;
		16'h37B8: out_word = 8'h31;
		16'h37B9: out_word = 8'h04;
		16'h37BA: out_word = 8'h31;
		16'h37BB: out_word = 8'h0F;
		16'h37BC: out_word = 8'hA1;
		16'h37BD: out_word = 8'h03;
		16'h37BE: out_word = 8'h86;
		16'h37BF: out_word = 8'h14;
		16'h37C0: out_word = 8'hE6;
		16'h37C1: out_word = 8'h5C;
		16'h37C2: out_word = 8'h1F;
		16'h37C3: out_word = 8'h0B;
		16'h37C4: out_word = 8'hA3;
		16'h37C5: out_word = 8'h8F;
		16'h37C6: out_word = 8'h38;
		16'h37C7: out_word = 8'hEE;
		16'h37C8: out_word = 8'hE9;
		16'h37C9: out_word = 8'h15;
		16'h37CA: out_word = 8'h63;
		16'h37CB: out_word = 8'hBB;
		16'h37CC: out_word = 8'h23;
		16'h37CD: out_word = 8'hEE;
		16'h37CE: out_word = 8'h92;
		16'h37CF: out_word = 8'h0D;
		16'h37D0: out_word = 8'hCD;
		16'h37D1: out_word = 8'hED;
		16'h37D2: out_word = 8'hF1;
		16'h37D3: out_word = 8'h23;
		16'h37D4: out_word = 8'h5D;
		16'h37D5: out_word = 8'h1B;
		16'h37D6: out_word = 8'hEA;
		16'h37D7: out_word = 8'h04;
		16'h37D8: out_word = 8'h38;
		16'h37D9: out_word = 8'hC9;
		16'h37DA: out_word = 8'hEF;
		16'h37DB: out_word = 8'h31;
		16'h37DC: out_word = 8'h1F;
		16'h37DD: out_word = 8'h01;
		16'h37DE: out_word = 8'h20;
		16'h37DF: out_word = 8'h05;
		16'h37E0: out_word = 8'h38;
		16'h37E1: out_word = 8'hC9;
		16'h37E2: out_word = 8'hCD;
		16'h37E3: out_word = 8'h97;
		16'h37E4: out_word = 8'h32;
		16'h37E5: out_word = 8'h7E;
		16'h37E6: out_word = 8'hFE;
		16'h37E7: out_word = 8'h81;
		16'h37E8: out_word = 8'h38;
		16'h37E9: out_word = 8'h0E;
		16'h37EA: out_word = 8'hEF;
		16'h37EB: out_word = 8'hA1;
		16'h37EC: out_word = 8'h1B;
		16'h37ED: out_word = 8'h01;
		16'h37EE: out_word = 8'h05;
		16'h37EF: out_word = 8'h31;
		16'h37F0: out_word = 8'h36;
		16'h37F1: out_word = 8'hA3;
		16'h37F2: out_word = 8'h01;
		16'h37F3: out_word = 8'h00;
		16'h37F4: out_word = 8'h06;
		16'h37F5: out_word = 8'h1B;
		16'h37F6: out_word = 8'h33;
		16'h37F7: out_word = 8'h03;
		16'h37F8: out_word = 8'hEF;
		16'h37F9: out_word = 8'hA0;
		16'h37FA: out_word = 8'h01;
		16'h37FB: out_word = 8'h31;
		16'h37FC: out_word = 8'h31;
		16'h37FD: out_word = 8'h04;
		16'h37FE: out_word = 8'h31;
		16'h37FF: out_word = 8'h0F;
		16'h3800: out_word = 8'hA1;
		16'h3801: out_word = 8'h03;
		16'h3802: out_word = 8'h8C;
		16'h3803: out_word = 8'h10;
		16'h3804: out_word = 8'hB2;
		16'h3805: out_word = 8'h13;
		16'h3806: out_word = 8'h0E;
		16'h3807: out_word = 8'h55;
		16'h3808: out_word = 8'hE4;
		16'h3809: out_word = 8'h8D;
		16'h380A: out_word = 8'h58;
		16'h380B: out_word = 8'h39;
		16'h380C: out_word = 8'hBC;
		16'h380D: out_word = 8'h5B;
		16'h380E: out_word = 8'h98;
		16'h380F: out_word = 8'hFD;
		16'h3810: out_word = 8'h9E;
		16'h3811: out_word = 8'h00;
		16'h3812: out_word = 8'h36;
		16'h3813: out_word = 8'h75;
		16'h3814: out_word = 8'hA0;
		16'h3815: out_word = 8'hDB;
		16'h3816: out_word = 8'hE8;
		16'h3817: out_word = 8'hB4;
		16'h3818: out_word = 8'h63;
		16'h3819: out_word = 8'h42;
		16'h381A: out_word = 8'hC4;
		16'h381B: out_word = 8'hE6;
		16'h381C: out_word = 8'hB5;
		16'h381D: out_word = 8'h09;
		16'h381E: out_word = 8'h36;
		16'h381F: out_word = 8'hBE;
		16'h3820: out_word = 8'hE9;
		16'h3821: out_word = 8'h36;
		16'h3822: out_word = 8'h73;
		16'h3823: out_word = 8'h1B;
		16'h3824: out_word = 8'h5D;
		16'h3825: out_word = 8'hEC;
		16'h3826: out_word = 8'hD8;
		16'h3827: out_word = 8'hDE;
		16'h3828: out_word = 8'h63;
		16'h3829: out_word = 8'hBE;
		16'h382A: out_word = 8'hF0;
		16'h382B: out_word = 8'h61;
		16'h382C: out_word = 8'hA1;
		16'h382D: out_word = 8'hB3;
		16'h382E: out_word = 8'h0C;
		16'h382F: out_word = 8'h04;
		16'h3830: out_word = 8'h0F;
		16'h3831: out_word = 8'h38;
		16'h3832: out_word = 8'hC9;
		16'h3833: out_word = 8'hEF;
		16'h3834: out_word = 8'h31;
		16'h3835: out_word = 8'h31;
		16'h3836: out_word = 8'h04;
		16'h3837: out_word = 8'hA1;
		16'h3838: out_word = 8'h03;
		16'h3839: out_word = 8'h1B;
		16'h383A: out_word = 8'h28;
		16'h383B: out_word = 8'hA1;
		16'h383C: out_word = 8'h0F;
		16'h383D: out_word = 8'h05;
		16'h383E: out_word = 8'h24;
		16'h383F: out_word = 8'h31;
		16'h3840: out_word = 8'h0F;
		16'h3841: out_word = 8'h38;
		16'h3842: out_word = 8'hC9;
		16'h3843: out_word = 8'hEF;
		16'h3844: out_word = 8'h22;
		16'h3845: out_word = 8'hA3;
		16'h3846: out_word = 8'h03;
		16'h3847: out_word = 8'h1B;
		16'h3848: out_word = 8'h38;
		16'h3849: out_word = 8'hC9;
		16'h384A: out_word = 8'hEF;
		16'h384B: out_word = 8'h31;
		16'h384C: out_word = 8'h30;
		16'h384D: out_word = 8'h00;
		16'h384E: out_word = 8'h1E;
		16'h384F: out_word = 8'hA2;
		16'h3850: out_word = 8'h38;
		16'h3851: out_word = 8'hEF;
		16'h3852: out_word = 8'h01;
		16'h3853: out_word = 8'h31;
		16'h3854: out_word = 8'h30;
		16'h3855: out_word = 8'h00;
		16'h3856: out_word = 8'h07;
		16'h3857: out_word = 8'h25;
		16'h3858: out_word = 8'h04;
		16'h3859: out_word = 8'h38;
		16'h385A: out_word = 8'hC3;
		16'h385B: out_word = 8'hC4;
		16'h385C: out_word = 8'h36;
		16'h385D: out_word = 8'h02;
		16'h385E: out_word = 8'h31;
		16'h385F: out_word = 8'h30;
		16'h3860: out_word = 8'h00;
		16'h3861: out_word = 8'h09;
		16'h3862: out_word = 8'hA0;
		16'h3863: out_word = 8'h01;
		16'h3864: out_word = 8'h37;
		16'h3865: out_word = 8'h00;
		16'h3866: out_word = 8'h06;
		16'h3867: out_word = 8'hA1;
		16'h3868: out_word = 8'h01;
		16'h3869: out_word = 8'h05;
		16'h386A: out_word = 8'h02;
		16'h386B: out_word = 8'hA1;
		16'h386C: out_word = 8'h38;
		16'h386D: out_word = 8'hC9;
		16'h386E: out_word = 8'hDD;
		16'h386F: out_word = 8'hE5;
		16'h3870: out_word = 8'hFD;
		16'h3871: out_word = 8'hCB;
		16'h3872: out_word = 8'h01;
		16'h3873: out_word = 8'h66;
		16'h3874: out_word = 8'h28;
		16'h3875: out_word = 8'h03;
		16'h3876: out_word = 8'hCD;
		16'h3877: out_word = 8'h42;
		16'h3878: out_word = 8'h3A;
		16'h3879: out_word = 8'hCD;
		16'h387A: out_word = 8'hBF;
		16'h387B: out_word = 8'h02;
		16'h387C: out_word = 8'hDD;
		16'h387D: out_word = 8'hE1;
		16'h387E: out_word = 8'hC9;
		16'h387F: out_word = 8'h0E;
		16'h3880: out_word = 8'hFD;
		16'h3881: out_word = 8'h16;
		16'h3882: out_word = 8'hFF;
		16'h3883: out_word = 8'h1E;
		16'h3884: out_word = 8'hBF;
		16'h3885: out_word = 8'h42;
		16'h3886: out_word = 8'h3E;
		16'h3887: out_word = 8'h07;
		16'h3888: out_word = 8'hED;
		16'h3889: out_word = 8'h79;
		16'h388A: out_word = 8'hED;
		16'h388B: out_word = 8'h60;
		16'h388C: out_word = 8'h3E;
		16'h388D: out_word = 8'h0E;
		16'h388E: out_word = 8'hED;
		16'h388F: out_word = 8'h79;
		16'h3890: out_word = 8'hED;
		16'h3891: out_word = 8'h78;
		16'h3892: out_word = 8'hF6;
		16'h3893: out_word = 8'hF0;
		16'h3894: out_word = 8'h6F;
		16'h3895: out_word = 8'hC9;
		16'h3896: out_word = 8'h42;
		16'h3897: out_word = 8'h3E;
		16'h3898: out_word = 8'h0E;
		16'h3899: out_word = 8'hED;
		16'h389A: out_word = 8'h79;
		16'h389B: out_word = 8'h43;
		16'h389C: out_word = 8'hED;
		16'h389D: out_word = 8'h69;
		16'h389E: out_word = 8'hC9;
		16'h389F: out_word = 8'h42;
		16'h38A0: out_word = 8'h3E;
		16'h38A1: out_word = 8'h0E;
		16'h38A2: out_word = 8'hED;
		16'h38A3: out_word = 8'h79;
		16'h38A4: out_word = 8'hED;
		16'h38A5: out_word = 8'h78;
		16'h38A6: out_word = 8'hC9;
		16'h38A7: out_word = 8'h7D;
		16'h38A8: out_word = 8'hE6;
		16'h38A9: out_word = 8'hFE;
		16'h38AA: out_word = 8'h6F;
		16'h38AB: out_word = 8'h18;
		16'h38AC: out_word = 8'hE9;
		16'h38AD: out_word = 8'h7D;
		16'h38AE: out_word = 8'hF6;
		16'h38AF: out_word = 8'h01;
		16'h38B0: out_word = 8'h6F;
		16'h38B1: out_word = 8'h18;
		16'h38B2: out_word = 8'hE3;
		16'h38B3: out_word = 8'h10;
		16'h38B4: out_word = 8'hFE;
		16'h38B5: out_word = 8'hC9;
		16'h38B6: out_word = 8'hC5;
		16'h38B7: out_word = 8'h06;
		16'h38B8: out_word = 8'h10;
		16'h38B9: out_word = 8'hCD;
		16'h38BA: out_word = 8'hB3;
		16'h38BB: out_word = 8'h38;
		16'h38BC: out_word = 8'hC1;
		16'h38BD: out_word = 8'h10;
		16'h38BE: out_word = 8'hF7;
		16'h38BF: out_word = 8'hC9;
		16'h38C0: out_word = 8'hC5;
		16'h38C1: out_word = 8'hCD;
		16'h38C2: out_word = 8'h9F;
		16'h38C3: out_word = 8'h38;
		16'h38C4: out_word = 8'hC1;
		16'h38C5: out_word = 8'hE6;
		16'h38C6: out_word = 8'h20;
		16'h38C7: out_word = 8'h28;
		16'h38C8: out_word = 8'h02;
		16'h38C9: out_word = 8'h10;
		16'h38CA: out_word = 8'hF5;
		16'h38CB: out_word = 8'hC9;
		16'h38CC: out_word = 8'hC5;
		16'h38CD: out_word = 8'hCD;
		16'h38CE: out_word = 8'h9F;
		16'h38CF: out_word = 8'h38;
		16'h38D0: out_word = 8'hC1;
		16'h38D1: out_word = 8'hE6;
		16'h38D2: out_word = 8'h20;
		16'h38D3: out_word = 8'h20;
		16'h38D4: out_word = 8'h02;
		16'h38D5: out_word = 8'h10;
		16'h38D6: out_word = 8'hF5;
		16'h38D7: out_word = 8'hC9;
		16'h38D8: out_word = 8'hCD;
		16'h38D9: out_word = 8'h7F;
		16'h38DA: out_word = 8'h38;
		16'h38DB: out_word = 8'h06;
		16'h38DC: out_word = 8'h01;
		16'h38DD: out_word = 8'h18;
		16'h38DE: out_word = 8'h05;
		16'h38DF: out_word = 8'hCD;
		16'h38E0: out_word = 8'h7F;
		16'h38E1: out_word = 8'h38;
		16'h38E2: out_word = 8'h06;
		16'h38E3: out_word = 8'h04;
		16'h38E4: out_word = 8'hC5;
		16'h38E5: out_word = 8'hCD;
		16'h38E6: out_word = 8'h9F;
		16'h38E7: out_word = 8'h38;
		16'h38E8: out_word = 8'hC1;
		16'h38E9: out_word = 8'hE6;
		16'h38EA: out_word = 8'h20;
		16'h38EB: out_word = 8'h28;
		16'h38EC: out_word = 8'h40;
		16'h38ED: out_word = 8'hAF;
		16'h38EE: out_word = 8'hC5;
		16'h38EF: out_word = 8'hF5;
		16'h38F0: out_word = 8'hCD;
		16'h38F1: out_word = 8'hAD;
		16'h38F2: out_word = 8'h38;
		16'h38F3: out_word = 8'h06;
		16'h38F4: out_word = 8'hA3;
		16'h38F5: out_word = 8'hCD;
		16'h38F6: out_word = 8'hC0;
		16'h38F7: out_word = 8'h38;
		16'h38F8: out_word = 8'h20;
		16'h38F9: out_word = 8'h31;
		16'h38FA: out_word = 8'hCD;
		16'h38FB: out_word = 8'hA7;
		16'h38FC: out_word = 8'h38;
		16'h38FD: out_word = 8'h18;
		16'h38FE: out_word = 8'h02;
		16'h38FF: out_word = 8'hFF;
		16'h3900: out_word = 8'hFF;
		16'h3901: out_word = 8'h06;
		16'h3902: out_word = 8'h2B;
		16'h3903: out_word = 8'hCD;
		16'h3904: out_word = 8'hB3;
		16'h3905: out_word = 8'h38;
		16'h3906: out_word = 8'hCD;
		16'h3907: out_word = 8'h9F;
		16'h3908: out_word = 8'h38;
		16'h3909: out_word = 8'hCB;
		16'h390A: out_word = 8'h6F;
		16'h390B: out_word = 8'h28;
		16'h390C: out_word = 8'h04;
		16'h390D: out_word = 8'hF1;
		16'h390E: out_word = 8'h37;
		16'h390F: out_word = 8'h18;
		16'h3910: out_word = 8'h03;
		16'h3911: out_word = 8'hF1;
		16'h3912: out_word = 8'h37;
		16'h3913: out_word = 8'h3F;
		16'h3914: out_word = 8'h1F;
		16'h3915: out_word = 8'hF5;
		16'h3916: out_word = 8'hCD;
		16'h3917: out_word = 8'hAD;
		16'h3918: out_word = 8'h38;
		16'h3919: out_word = 8'h06;
		16'h391A: out_word = 8'h26;
		16'h391B: out_word = 8'hCD;
		16'h391C: out_word = 8'hB3;
		16'h391D: out_word = 8'h38;
		16'h391E: out_word = 8'hCD;
		16'h391F: out_word = 8'hA7;
		16'h3920: out_word = 8'h38;
		16'h3921: out_word = 8'h06;
		16'h3922: out_word = 8'h23;
		16'h3923: out_word = 8'hCD;
		16'h3924: out_word = 8'hB3;
		16'h3925: out_word = 8'h38;
		16'h3926: out_word = 8'hF1;
		16'h3927: out_word = 8'hC1;
		16'h3928: out_word = 8'h10;
		16'h3929: out_word = 8'hC4;
		16'h392A: out_word = 8'hC9;
		16'h392B: out_word = 8'hF1;
		16'h392C: out_word = 8'hC1;
		16'h392D: out_word = 8'hCD;
		16'h392E: out_word = 8'hAD;
		16'h392F: out_word = 8'h38;
		16'h3930: out_word = 8'hAF;
		16'h3931: out_word = 8'h32;
		16'h3932: out_word = 8'h88;
		16'h3933: out_word = 8'h5B;
		16'h3934: out_word = 8'h3C;
		16'h3935: out_word = 8'h37;
		16'h3936: out_word = 8'h3F;
		16'h3937: out_word = 8'hC9;
		16'h3938: out_word = 8'hCD;
		16'h3939: out_word = 8'h7F;
		16'h393A: out_word = 8'h38;
		16'h393B: out_word = 8'h3A;
		16'h393C: out_word = 8'h88;
		16'h393D: out_word = 8'h5B;
		16'h393E: out_word = 8'hE6;
		16'h393F: out_word = 8'h80;
		16'h3940: out_word = 8'h20;
		16'h3941: out_word = 8'h57;
		16'h3942: out_word = 8'hCD;
		16'h3943: out_word = 8'h9F;
		16'h3944: out_word = 8'h38;
		16'h3945: out_word = 8'hE6;
		16'h3946: out_word = 8'h20;
		16'h3947: out_word = 8'h28;
		16'h3948: out_word = 8'hE4;
		16'h3949: out_word = 8'h3A;
		16'h394A: out_word = 8'h88;
		16'h394B: out_word = 8'h5B;
		16'h394C: out_word = 8'hA7;
		16'h394D: out_word = 8'h20;
		16'h394E: out_word = 8'h0B;
		16'h394F: out_word = 8'h3C;
		16'h3950: out_word = 8'h32;
		16'h3951: out_word = 8'h88;
		16'h3952: out_word = 8'h5B;
		16'h3953: out_word = 8'h3E;
		16'h3954: out_word = 8'h4C;
		16'h3955: out_word = 8'h32;
		16'h3956: out_word = 8'h89;
		16'h3957: out_word = 8'h5B;
		16'h3958: out_word = 8'h18;
		16'h3959: out_word = 8'h42;
		16'h395A: out_word = 8'h3A;
		16'h395B: out_word = 8'h89;
		16'h395C: out_word = 8'h5B;
		16'h395D: out_word = 8'h3D;
		16'h395E: out_word = 8'h32;
		16'h395F: out_word = 8'h89;
		16'h3960: out_word = 8'h5B;
		16'h3961: out_word = 8'h20;
		16'h3962: out_word = 8'h39;
		16'h3963: out_word = 8'hAF;
		16'h3964: out_word = 8'h32;
		16'h3965: out_word = 8'h88;
		16'h3966: out_word = 8'h5B;
		16'h3967: out_word = 8'h32;
		16'h3968: out_word = 8'h89;
		16'h3969: out_word = 8'h5B;
		16'h396A: out_word = 8'h32;
		16'h396B: out_word = 8'h8A;
		16'h396C: out_word = 8'h5B;
		16'h396D: out_word = 8'hCD;
		16'h396E: out_word = 8'hA7;
		16'h396F: out_word = 8'h38;
		16'h3970: out_word = 8'h06;
		16'h3971: out_word = 8'h21;
		16'h3972: out_word = 8'hCD;
		16'h3973: out_word = 8'hC0;
		16'h3974: out_word = 8'h38;
		16'h3975: out_word = 8'h20;
		16'h3976: out_word = 8'hB6;
		16'h3977: out_word = 8'hCD;
		16'h3978: out_word = 8'hAD;
		16'h3979: out_word = 8'h38;
		16'h397A: out_word = 8'h06;
		16'h397B: out_word = 8'h24;
		16'h397C: out_word = 8'hCD;
		16'h397D: out_word = 8'hCC;
		16'h397E: out_word = 8'h38;
		16'h397F: out_word = 8'h28;
		16'h3980: out_word = 8'hAC;
		16'h3981: out_word = 8'hCD;
		16'h3982: out_word = 8'hA7;
		16'h3983: out_word = 8'h38;
		16'h3984: out_word = 8'h06;
		16'h3985: out_word = 8'h0F;
		16'h3986: out_word = 8'hCD;
		16'h3987: out_word = 8'hB6;
		16'h3988: out_word = 8'h38;
		16'h3989: out_word = 8'hCD;
		16'h398A: out_word = 8'hDF;
		16'h398B: out_word = 8'h38;
		16'h398C: out_word = 8'h20;
		16'h398D: out_word = 8'h9F;
		16'h398E: out_word = 8'hCB;
		16'h398F: out_word = 8'hFF;
		16'h3990: out_word = 8'hE6;
		16'h3991: out_word = 8'hF0;
		16'h3992: out_word = 8'h32;
		16'h3993: out_word = 8'h88;
		16'h3994: out_word = 8'h5B;
		16'h3995: out_word = 8'hAF;
		16'h3996: out_word = 8'hCB;
		16'h3997: out_word = 8'h3F;
		16'h3998: out_word = 8'hC9;
		16'h3999: out_word = 8'hAF;
		16'h399A: out_word = 8'h37;
		16'h399B: out_word = 8'hC9;
		16'h399C: out_word = 8'hAF;
		16'h399D: out_word = 8'h3C;
		16'h399E: out_word = 8'h37;
		16'h399F: out_word = 8'hC9;
		16'h39A0: out_word = 8'hCD;
		16'h39A1: out_word = 8'h38;
		16'h39A2: out_word = 8'h39;
		16'h39A3: out_word = 8'h3A;
		16'h39A4: out_word = 8'h88;
		16'h39A5: out_word = 8'h5B;
		16'h39A6: out_word = 8'h2F;
		16'h39A7: out_word = 8'hE6;
		16'h39A8: out_word = 8'hC0;
		16'h39A9: out_word = 8'hC0;
		16'h39AA: out_word = 8'hDD;
		16'h39AB: out_word = 8'h21;
		16'h39AC: out_word = 8'h8A;
		16'h39AD: out_word = 8'h5B;
		16'h39AE: out_word = 8'h06;
		16'h39AF: out_word = 8'h05;
		16'h39B0: out_word = 8'hC5;
		16'h39B1: out_word = 8'hCD;
		16'h39B2: out_word = 8'hD8;
		16'h39B3: out_word = 8'h38;
		16'h39B4: out_word = 8'hC2;
		16'h39B5: out_word = 8'h3A;
		16'h39B6: out_word = 8'h3A;
		16'h39B7: out_word = 8'hCB;
		16'h39B8: out_word = 8'h7F;
		16'h39B9: out_word = 8'h28;
		16'h39BA: out_word = 8'h21;
		16'h39BB: out_word = 8'hCD;
		16'h39BC: out_word = 8'hDF;
		16'h39BD: out_word = 8'h38;
		16'h39BE: out_word = 8'h20;
		16'h39BF: out_word = 8'h7A;
		16'h39C0: out_word = 8'hC1;
		16'h39C1: out_word = 8'hC5;
		16'h39C2: out_word = 8'h4F;
		16'h39C3: out_word = 8'hDD;
		16'h39C4: out_word = 8'h7E;
		16'h39C5: out_word = 8'h00;
		16'h39C6: out_word = 8'hCB;
		16'h39C7: out_word = 8'h40;
		16'h39C8: out_word = 8'h28;
		16'h39C9: out_word = 8'h0C;
		16'h39CA: out_word = 8'hCB;
		16'h39CB: out_word = 8'h39;
		16'h39CC: out_word = 8'hCB;
		16'h39CD: out_word = 8'h39;
		16'h39CE: out_word = 8'hCB;
		16'h39CF: out_word = 8'h39;
		16'h39D0: out_word = 8'hCB;
		16'h39D1: out_word = 8'h39;
		16'h39D2: out_word = 8'hE6;
		16'h39D3: out_word = 8'hF0;
		16'h39D4: out_word = 8'h18;
		16'h39D5: out_word = 8'h02;
		16'h39D6: out_word = 8'hE6;
		16'h39D7: out_word = 8'h0F;
		16'h39D8: out_word = 8'hB1;
		16'h39D9: out_word = 8'hDD;
		16'h39DA: out_word = 8'h77;
		16'h39DB: out_word = 8'h00;
		16'h39DC: out_word = 8'hC1;
		16'h39DD: out_word = 8'hCB;
		16'h39DE: out_word = 8'h40;
		16'h39DF: out_word = 8'h20;
		16'h39E0: out_word = 8'h02;
		16'h39E1: out_word = 8'hDD;
		16'h39E2: out_word = 8'h2B;
		16'h39E3: out_word = 8'h10;
		16'h39E4: out_word = 8'hCB;
		16'h39E5: out_word = 8'h1E;
		16'h39E6: out_word = 8'h80;
		16'h39E7: out_word = 8'hDD;
		16'h39E8: out_word = 8'h21;
		16'h39E9: out_word = 8'h88;
		16'h39EA: out_word = 8'h5B;
		16'h39EB: out_word = 8'h21;
		16'h39EC: out_word = 8'h3F;
		16'h39ED: out_word = 8'h3A;
		16'h39EE: out_word = 8'h06;
		16'h39EF: out_word = 8'h03;
		16'h39F0: out_word = 8'hDD;
		16'h39F1: out_word = 8'h7E;
		16'h39F2: out_word = 8'h00;
		16'h39F3: out_word = 8'hA6;
		16'h39F4: out_word = 8'h28;
		16'h39F5: out_word = 8'h21;
		16'h39F6: out_word = 8'hCB;
		16'h39F7: out_word = 8'h7B;
		16'h39F8: out_word = 8'h28;
		16'h39F9: out_word = 8'h42;
		16'h39FA: out_word = 8'hC5;
		16'h39FB: out_word = 8'hF5;
		16'h39FC: out_word = 8'h78;
		16'h39FD: out_word = 8'h18;
		16'h39FE: out_word = 8'h02;
		16'h39FF: out_word = 8'hFF;
		16'h3A00: out_word = 8'hFF;
		16'h3A01: out_word = 8'h3D;
		16'h3A02: out_word = 8'hCB;
		16'h3A03: out_word = 8'h27;
		16'h3A04: out_word = 8'hCB;
		16'h3A05: out_word = 8'h27;
		16'h3A06: out_word = 8'hCB;
		16'h3A07: out_word = 8'h27;
		16'h3A08: out_word = 8'hF6;
		16'h3A09: out_word = 8'h07;
		16'h3A0A: out_word = 8'h47;
		16'h3A0B: out_word = 8'hF1;
		16'h3A0C: out_word = 8'hCB;
		16'h3A0D: out_word = 8'h27;
		16'h3A0E: out_word = 8'hDA;
		16'h3A0F: out_word = 8'h13;
		16'h3A10: out_word = 8'h3A;
		16'h3A11: out_word = 8'h10;
		16'h3A12: out_word = 8'hF9;
		16'h3A13: out_word = 8'h58;
		16'h3A14: out_word = 8'hC1;
		16'h3A15: out_word = 8'h20;
		16'h3A16: out_word = 8'h25;
		16'h3A17: out_word = 8'hDD;
		16'h3A18: out_word = 8'h23;
		16'h3A19: out_word = 8'h23;
		16'h3A1A: out_word = 8'h10;
		16'h3A1B: out_word = 8'hD4;
		16'h3A1C: out_word = 8'hCB;
		16'h3A1D: out_word = 8'h7B;
		16'h3A1E: out_word = 8'h20;
		16'h3A1F: out_word = 8'h07;
		16'h3A20: out_word = 8'h7B;
		16'h3A21: out_word = 8'hE6;
		16'h3A22: out_word = 8'hFC;
		16'h3A23: out_word = 8'h28;
		16'h3A24: out_word = 8'h02;
		16'h3A25: out_word = 8'h1D;
		16'h3A26: out_word = 8'h1D;
		16'h3A27: out_word = 8'h3A;
		16'h3A28: out_word = 8'h8A;
		16'h3A29: out_word = 8'h5B;
		16'h3A2A: out_word = 8'hE6;
		16'h3A2B: out_word = 8'h08;
		16'h3A2C: out_word = 8'h28;
		16'h3A2D: out_word = 8'h06;
		16'h3A2E: out_word = 8'h7B;
		16'h3A2F: out_word = 8'hE6;
		16'h3A30: out_word = 8'h7F;
		16'h3A31: out_word = 8'hC6;
		16'h3A32: out_word = 8'h12;
		16'h3A33: out_word = 8'h5F;
		16'h3A34: out_word = 8'h7B;
		16'h3A35: out_word = 8'hC6;
		16'h3A36: out_word = 8'h5A;
		16'h3A37: out_word = 8'h5F;
		16'h3A38: out_word = 8'hAF;
		16'h3A39: out_word = 8'hC9;
		16'h3A3A: out_word = 8'hC1;
		16'h3A3B: out_word = 8'hC9;
		16'h3A3C: out_word = 8'hAF;
		16'h3A3D: out_word = 8'h3C;
		16'h3A3E: out_word = 8'hC9;
		16'h3A3F: out_word = 8'h0F;
		16'h3A40: out_word = 8'hFF;
		16'h3A41: out_word = 8'hF2;
		16'h3A42: out_word = 8'h1E;
		16'h3A43: out_word = 8'h80;
		16'h3A44: out_word = 8'h3A;
		16'h3A45: out_word = 8'h78;
		16'h3A46: out_word = 8'h5C;
		16'h3A47: out_word = 8'hE6;
		16'h3A48: out_word = 8'h01;
		16'h3A49: out_word = 8'h20;
		16'h3A4A: out_word = 8'h04;
		16'h3A4B: out_word = 8'hCD;
		16'h3A4C: out_word = 8'hA0;
		16'h3A4D: out_word = 8'h39;
		16'h3A4E: out_word = 8'hC0;
		16'h3A4F: out_word = 8'h21;
		16'h3A50: out_word = 8'h00;
		16'h3A51: out_word = 8'h5C;
		16'h3A52: out_word = 8'hCB;
		16'h3A53: out_word = 8'h7E;
		16'h3A54: out_word = 8'h20;
		16'h3A55: out_word = 8'h0C;
		16'h3A56: out_word = 8'h7E;
		16'h3A57: out_word = 8'hFE;
		16'h3A58: out_word = 8'h5B;
		16'h3A59: out_word = 8'h38;
		16'h3A5A: out_word = 8'h07;
		16'h3A5B: out_word = 8'h23;
		16'h3A5C: out_word = 8'h35;
		16'h3A5D: out_word = 8'h2B;
		16'h3A5E: out_word = 8'h20;
		16'h3A5F: out_word = 8'h02;
		16'h3A60: out_word = 8'h36;
		16'h3A61: out_word = 8'hFF;
		16'h3A62: out_word = 8'h7D;
		16'h3A63: out_word = 8'h21;
		16'h3A64: out_word = 8'h04;
		16'h3A65: out_word = 8'h5C;
		16'h3A66: out_word = 8'hBD;
		16'h3A67: out_word = 8'h20;
		16'h3A68: out_word = 8'hE9;
		16'h3A69: out_word = 8'hCD;
		16'h3A6A: out_word = 8'hAE;
		16'h3A6B: out_word = 8'h3A;
		16'h3A6C: out_word = 8'hC0;
		16'h3A6D: out_word = 8'h7B;
		16'h3A6E: out_word = 8'h21;
		16'h3A6F: out_word = 8'h00;
		16'h3A70: out_word = 8'h5C;
		16'h3A71: out_word = 8'hBE;
		16'h3A72: out_word = 8'h28;
		16'h3A73: out_word = 8'h2A;
		16'h3A74: out_word = 8'hEB;
		16'h3A75: out_word = 8'h21;
		16'h3A76: out_word = 8'h04;
		16'h3A77: out_word = 8'h5C;
		16'h3A78: out_word = 8'hBE;
		16'h3A79: out_word = 8'h28;
		16'h3A7A: out_word = 8'h23;
		16'h3A7B: out_word = 8'hCB;
		16'h3A7C: out_word = 8'h7E;
		16'h3A7D: out_word = 8'h20;
		16'h3A7E: out_word = 8'h04;
		16'h3A7F: out_word = 8'hEB;
		16'h3A80: out_word = 8'hCB;
		16'h3A81: out_word = 8'h7E;
		16'h3A82: out_word = 8'hC8;
		16'h3A83: out_word = 8'h5F;
		16'h3A84: out_word = 8'h77;
		16'h3A85: out_word = 8'h23;
		16'h3A86: out_word = 8'h36;
		16'h3A87: out_word = 8'h0A;
		16'h3A88: out_word = 8'h23;
		16'h3A89: out_word = 8'h3A;
		16'h3A8A: out_word = 8'h09;
		16'h3A8B: out_word = 8'h5C;
		16'h3A8C: out_word = 8'hCB;
		16'h3A8D: out_word = 8'h3F;
		16'h3A8E: out_word = 8'h77;
		16'h3A8F: out_word = 8'h23;
		16'h3A90: out_word = 8'hCD;
		16'h3A91: out_word = 8'hD7;
		16'h3A92: out_word = 8'h3A;
		16'h3A93: out_word = 8'h73;
		16'h3A94: out_word = 8'h7B;
		16'h3A95: out_word = 8'h32;
		16'h3A96: out_word = 8'h08;
		16'h3A97: out_word = 8'h5C;
		16'h3A98: out_word = 8'h21;
		16'h3A99: out_word = 8'h3B;
		16'h3A9A: out_word = 8'h5C;
		16'h3A9B: out_word = 8'hCB;
		16'h3A9C: out_word = 8'hEE;
		16'h3A9D: out_word = 8'hC9;
		16'h3A9E: out_word = 8'h23;
		16'h3A9F: out_word = 8'h36;
		16'h3AA0: out_word = 8'h0A;
		16'h3AA1: out_word = 8'h23;
		16'h3AA2: out_word = 8'h35;
		16'h3AA3: out_word = 8'hC0;
		16'h3AA4: out_word = 8'h3A;
		16'h3AA5: out_word = 8'h0A;
		16'h3AA6: out_word = 8'h5C;
		16'h3AA7: out_word = 8'hCB;
		16'h3AA8: out_word = 8'h3F;
		16'h3AA9: out_word = 8'h77;
		16'h3AAA: out_word = 8'h23;
		16'h3AAB: out_word = 8'h5E;
		16'h3AAC: out_word = 8'h18;
		16'h3AAD: out_word = 8'hE6;
		16'h3AAE: out_word = 8'h7B;
		16'h3AAF: out_word = 8'h21;
		16'h3AB0: out_word = 8'h66;
		16'h3AB1: out_word = 8'h5B;
		16'h3AB2: out_word = 8'hCB;
		16'h3AB3: out_word = 8'h46;
		16'h3AB4: out_word = 8'h28;
		16'h3AB5: out_word = 8'h06;
		16'h3AB6: out_word = 8'hFE;
		16'h3AB7: out_word = 8'h6D;
		16'h3AB8: out_word = 8'h30;
		16'h3AB9: out_word = 8'h1A;
		16'h3ABA: out_word = 8'hAF;
		16'h3ABB: out_word = 8'hC9;
		16'h3ABC: out_word = 8'hFE;
		16'h3ABD: out_word = 8'h80;
		16'h3ABE: out_word = 8'h30;
		16'h3ABF: out_word = 8'h14;
		16'h3AC0: out_word = 8'hFE;
		16'h3AC1: out_word = 8'h6C;
		16'h3AC2: out_word = 8'h20;
		16'h3AC3: out_word = 8'hF6;
		16'h3AC4: out_word = 8'h00;
		16'h3AC5: out_word = 8'h00;
		16'h3AC6: out_word = 8'h00;
		16'h3AC7: out_word = 8'h00;
		16'h3AC8: out_word = 8'h00;
		16'h3AC9: out_word = 8'h00;
		16'h3ACA: out_word = 8'h00;
		16'h3ACB: out_word = 8'h00;
		16'h3ACC: out_word = 8'h00;
		16'h3ACD: out_word = 8'h00;
		16'h3ACE: out_word = 8'h00;
		16'h3ACF: out_word = 8'h00;
		16'h3AD0: out_word = 8'h00;
		16'h3AD1: out_word = 8'h00;
		16'h3AD2: out_word = 8'h00;
		16'h3AD3: out_word = 8'h00;
		16'h3AD4: out_word = 8'hAF;
		16'h3AD5: out_word = 8'h3C;
		16'h3AD6: out_word = 8'hC9;
		16'h3AD7: out_word = 8'hE5;
		16'h3AD8: out_word = 8'h7B;
		16'h3AD9: out_word = 8'hD6;
		16'h3ADA: out_word = 8'h5B;
		16'h3ADB: out_word = 8'h16;
		16'h3ADC: out_word = 8'h00;
		16'h3ADD: out_word = 8'h5F;
		16'h3ADE: out_word = 8'h21;
		16'h3ADF: out_word = 8'h66;
		16'h3AE0: out_word = 8'h5B;
		16'h3AE1: out_word = 8'hCB;
		16'h3AE2: out_word = 8'h46;
		16'h3AE3: out_word = 8'h28;
		16'h3AE4: out_word = 8'h05;
		16'h3AE5: out_word = 8'h21;
		16'h3AE6: out_word = 8'h13;
		16'h3AE7: out_word = 8'h3B;
		16'h3AE8: out_word = 8'h18;
		16'h3AE9: out_word = 8'h25;
		16'h3AEA: out_word = 8'h21;
		16'h3AEB: out_word = 8'h25;
		16'h3AEC: out_word = 8'h3B;
		16'h3AED: out_word = 8'hFE;
		16'h3AEE: out_word = 8'h11;
		16'h3AEF: out_word = 8'h38;
		16'h3AF0: out_word = 8'h1E;
		16'h3AF1: out_word = 8'h21;
		16'h3AF2: out_word = 8'h21;
		16'h3AF3: out_word = 8'h3B;
		16'h3AF4: out_word = 8'hFE;
		16'h3AF5: out_word = 8'h15;
		16'h3AF6: out_word = 8'h28;
		16'h3AF7: out_word = 8'h17;
		16'h3AF8: out_word = 8'hFE;
		16'h3AF9: out_word = 8'h16;
		16'h3AFA: out_word = 8'h28;
		16'h3AFB: out_word = 8'h13;
		16'h3AFC: out_word = 8'h18;
		16'h3AFD: out_word = 8'h03;
		16'h3AFE: out_word = 8'h00;
		16'h3AFF: out_word = 8'hFF;
		16'h3B00: out_word = 8'hFF;
		16'h3B01: out_word = 8'hFE;
		16'h3B02: out_word = 8'h17;
		16'h3B03: out_word = 8'h28;
		16'h3B04: out_word = 8'h0A;
		16'h3B05: out_word = 8'h21;
		16'h3B06: out_word = 8'h18;
		16'h3B07: out_word = 8'h3B;
		16'h3B08: out_word = 8'hFE;
		16'h3B09: out_word = 8'h21;
		16'h3B0A: out_word = 8'h30;
		16'h3B0B: out_word = 8'h03;
		16'h3B0C: out_word = 8'h21;
		16'h3B0D: out_word = 8'h13;
		16'h3B0E: out_word = 8'h3B;
		16'h3B0F: out_word = 8'h19;
		16'h3B10: out_word = 8'h5E;
		16'h3B11: out_word = 8'hE1;
		16'h3B12: out_word = 8'hC9;
		16'h3B13: out_word = 8'h2E;
		16'h3B14: out_word = 8'h0D;
		16'h3B15: out_word = 8'h33;
		16'h3B16: out_word = 8'h32;
		16'h3B17: out_word = 8'h31;
		16'h3B18: out_word = 8'h29;
		16'h3B19: out_word = 8'h28;
		16'h3B1A: out_word = 8'h2A;
		16'h3B1B: out_word = 8'h2F;
		16'h3B1C: out_word = 8'h2D;
		16'h3B1D: out_word = 8'h39;
		16'h3B1E: out_word = 8'h38;
		16'h3B1F: out_word = 8'h37;
		16'h3B20: out_word = 8'h2B;
		16'h3B21: out_word = 8'h36;
		16'h3B22: out_word = 8'h35;
		16'h3B23: out_word = 8'h34;
		16'h3B24: out_word = 8'h30;
		16'h3B25: out_word = 8'hA5;
		16'h3B26: out_word = 8'h0D;
		16'h3B27: out_word = 8'hA6;
		16'h3B28: out_word = 8'hA7;
		16'h3B29: out_word = 8'hA8;
		16'h3B2A: out_word = 8'hA9;
		16'h3B2B: out_word = 8'hAA;
		16'h3B2C: out_word = 8'h0B;
		16'h3B2D: out_word = 8'h0C;
		16'h3B2E: out_word = 8'h07;
		16'h3B2F: out_word = 8'h09;
		16'h3B30: out_word = 8'h0A;
		16'h3B31: out_word = 8'h08;
		16'h3B32: out_word = 8'hAC;
		16'h3B33: out_word = 8'hAD;
		16'h3B34: out_word = 8'hAE;
		16'h3B35: out_word = 8'hAF;
		16'h3B36: out_word = 8'hB0;
		16'h3B37: out_word = 8'hB1;
		16'h3B38: out_word = 8'hB2;
		16'h3B39: out_word = 8'hB3;
		16'h3B3A: out_word = 8'hB4;
		16'h3B3B: out_word = 8'hFD;
		16'h3B3C: out_word = 8'hCB;
		16'h3B3D: out_word = 8'h01;
		16'h3B3E: out_word = 8'h66;
		16'h3B3F: out_word = 8'h20;
		16'h3B40: out_word = 8'h05;
		16'h3B41: out_word = 8'hAF;
		16'h3B42: out_word = 8'h11;
		16'h3B43: out_word = 8'h36;
		16'h3B44: out_word = 8'h15;
		16'h3B45: out_word = 8'hC9;
		16'h3B46: out_word = 8'h21;
		16'h3B47: out_word = 8'h0F;
		16'h3B48: out_word = 8'h01;
		16'h3B49: out_word = 8'hE3;
		16'h3B4A: out_word = 8'hC3;
		16'h3B4B: out_word = 8'h00;
		16'h3B4C: out_word = 8'h5B;
		16'h3B4D: out_word = 8'hFD;
		16'h3B4E: out_word = 8'hCB;
		16'h3B4F: out_word = 8'h01;
		16'h3B50: out_word = 8'h66;
		16'h3B51: out_word = 8'h20;
		16'h3B52: out_word = 8'h05;
		16'h3B53: out_word = 8'hFD;
		16'h3B54: out_word = 8'hCB;
		16'h3B55: out_word = 8'h0A;
		16'h3B56: out_word = 8'h7E;
		16'h3B57: out_word = 8'hC9;
		16'h3B58: out_word = 8'h21;
		16'h3B59: out_word = 8'h12;
		16'h3B5A: out_word = 8'h01;
		16'h3B5B: out_word = 8'h18;
		16'h3B5C: out_word = 8'hEC;
		16'h3B5D: out_word = 8'hFD;
		16'h3B5E: out_word = 8'hCB;
		16'h3B5F: out_word = 8'h01;
		16'h3B60: out_word = 8'h66;
		16'h3B61: out_word = 8'h20;
		16'h3B62: out_word = 8'h04;
		16'h3B63: out_word = 8'hDF;
		16'h3B64: out_word = 8'hFE;
		16'h3B65: out_word = 8'h0D;
		16'h3B66: out_word = 8'hC9;
		16'h3B67: out_word = 8'h21;
		16'h3B68: out_word = 8'h15;
		16'h3B69: out_word = 8'h01;
		16'h3B6A: out_word = 8'h18;
		16'h3B6B: out_word = 8'hDD;
		16'h3B6C: out_word = 8'hCD;
		16'h3B6D: out_word = 8'h8E;
		16'h3B6E: out_word = 8'h02;
		16'h3B6F: out_word = 8'h0E;
		16'h3B70: out_word = 8'h00;
		16'h3B71: out_word = 8'h20;
		16'h3B72: out_word = 8'h0D;
		16'h3B73: out_word = 8'hCD;
		16'h3B74: out_word = 8'h1E;
		16'h3B75: out_word = 8'h03;
		16'h3B76: out_word = 8'h30;
		16'h3B77: out_word = 8'h08;
		16'h3B78: out_word = 8'h15;
		16'h3B79: out_word = 8'h5F;
		16'h3B7A: out_word = 8'hCD;
		16'h3B7B: out_word = 8'h33;
		16'h3B7C: out_word = 8'h03;
		16'h3B7D: out_word = 8'hC3;
		16'h3B7E: out_word = 8'h57;
		16'h3B7F: out_word = 8'h26;
		16'h3B80: out_word = 8'hFD;
		16'h3B81: out_word = 8'hCB;
		16'h3B82: out_word = 8'h01;
		16'h3B83: out_word = 8'h66;
		16'h3B84: out_word = 8'hCA;
		16'h3B85: out_word = 8'h60;
		16'h3B86: out_word = 8'h26;
		16'h3B87: out_word = 8'hF3;
		16'h3B88: out_word = 8'hCD;
		16'h3B89: out_word = 8'hA0;
		16'h3B8A: out_word = 8'h39;
		16'h3B8B: out_word = 8'hFB;
		16'h3B8C: out_word = 8'h20;
		16'h3B8D: out_word = 8'h0C;
		16'h3B8E: out_word = 8'hCD;
		16'h3B8F: out_word = 8'hAE;
		16'h3B90: out_word = 8'h3A;
		16'h3B91: out_word = 8'h20;
		16'h3B92: out_word = 8'h07;
		16'h3B93: out_word = 8'hCD;
		16'h3B94: out_word = 8'hD7;
		16'h3B95: out_word = 8'h3A;
		16'h3B96: out_word = 8'h7B;
		16'h3B97: out_word = 8'hC3;
		16'h3B98: out_word = 8'h57;
		16'h3B99: out_word = 8'h26;
		16'h3B9A: out_word = 8'h0E;
		16'h3B9B: out_word = 8'h00;
		16'h3B9C: out_word = 8'hC3;
		16'h3B9D: out_word = 8'h60;
		16'h3B9E: out_word = 8'h26;
		16'h3B9F: out_word = 8'hFE;
		16'h3BA0: out_word = 8'hA3;
		16'h3BA1: out_word = 8'h28;
		16'h3BA2: out_word = 8'h0C;
		16'h3BA3: out_word = 8'hFE;
		16'h3BA4: out_word = 8'hA4;
		16'h3BA5: out_word = 8'h28;
		16'h3BA6: out_word = 8'h08;
		16'h3BA7: out_word = 8'hD6;
		16'h3BA8: out_word = 8'hA5;
		16'h3BA9: out_word = 8'hD2;
		16'h3BAA: out_word = 8'h5F;
		16'h3BAB: out_word = 8'h0B;
		16'h3BAC: out_word = 8'hC3;
		16'h3BAD: out_word = 8'h56;
		16'h3BAE: out_word = 8'h0B;
		16'h3BAF: out_word = 8'hFD;
		16'h3BB0: out_word = 8'hCB;
		16'h3BB1: out_word = 8'h01;
		16'h3BB2: out_word = 8'h66;
		16'h3BB3: out_word = 8'h28;
		16'h3BB4: out_word = 8'hF2;
		16'h3BB5: out_word = 8'h11;
		16'h3BB6: out_word = 8'hC9;
		16'h3BB7: out_word = 8'h3B;
		16'h3BB8: out_word = 8'hD5;
		16'h3BB9: out_word = 8'hD6;
		16'h3BBA: out_word = 8'hA3;
		16'h3BBB: out_word = 8'h11;
		16'h3BBC: out_word = 8'hD2;
		16'h3BBD: out_word = 8'h3B;
		16'h3BBE: out_word = 8'h28;
		16'h3BBF: out_word = 8'h03;
		16'h3BC0: out_word = 8'h11;
		16'h3BC1: out_word = 8'hDA;
		16'h3BC2: out_word = 8'h3B;
		16'h3BC3: out_word = 8'h3E;
		16'h3BC4: out_word = 8'h04;
		16'h3BC5: out_word = 8'hF5;
		16'h3BC6: out_word = 8'hC3;
		16'h3BC7: out_word = 8'h17;
		16'h3BC8: out_word = 8'h0C;
		16'h3BC9: out_word = 8'h37;
		16'h3BCA: out_word = 8'hFD;
		16'h3BCB: out_word = 8'hCB;
		16'h3BCC: out_word = 8'h01;
		16'h3BCD: out_word = 8'h4E;
		16'h3BCE: out_word = 8'hC0;
		16'h3BCF: out_word = 8'hC3;
		16'h3BD0: out_word = 8'h03;
		16'h3BD1: out_word = 8'h0B;
		16'h3BD2: out_word = 8'h53;
		16'h3BD3: out_word = 8'h50;
		16'h3BD4: out_word = 8'h45;
		16'h3BD5: out_word = 8'h43;
		16'h3BD6: out_word = 8'h54;
		16'h3BD7: out_word = 8'h52;
		16'h3BD8: out_word = 8'h55;
		16'h3BD9: out_word = 8'hCD;
		16'h3BDA: out_word = 8'h50;
		16'h3BDB: out_word = 8'h4C;
		16'h3BDC: out_word = 8'h41;
		16'h3BDD: out_word = 8'hD9;
		16'h3BDE: out_word = 8'hC3;
		16'h3BDF: out_word = 8'h01;
		16'h3BE0: out_word = 8'h3C;
		16'h3BE1: out_word = 8'h00;
		16'h3BE2: out_word = 8'h00;
		16'h3BE3: out_word = 8'h00;
		16'h3BE4: out_word = 8'h00;
		16'h3BE5: out_word = 8'h00;
		16'h3BE6: out_word = 8'h00;
		16'h3BE7: out_word = 8'h00;
		16'h3BE8: out_word = 8'h00;
		16'h3BE9: out_word = 8'h00;
		16'h3BEA: out_word = 8'h00;
		16'h3BEB: out_word = 8'h00;
		16'h3BEC: out_word = 8'h00;
		16'h3BED: out_word = 8'h00;
		16'h3BEE: out_word = 8'h00;
		16'h3BEF: out_word = 8'h00;
		16'h3BF0: out_word = 8'h00;
		16'h3BF1: out_word = 8'h00;
		16'h3BF2: out_word = 8'h00;
		16'h3BF3: out_word = 8'h00;
		16'h3BF4: out_word = 8'h00;
		16'h3BF5: out_word = 8'h00;
		16'h3BF6: out_word = 8'h00;
		16'h3BF7: out_word = 8'h00;
		16'h3BF8: out_word = 8'h00;
		16'h3BF9: out_word = 8'h00;
		16'h3BFA: out_word = 8'h00;
		16'h3BFB: out_word = 8'h00;
		16'h3BFC: out_word = 8'h00;
		16'h3BFD: out_word = 8'h00;
		16'h3BFE: out_word = 8'h00;
		16'h3BFF: out_word = 8'hFF;
		16'h3C00: out_word = 8'hFF;
		16'h3C01: out_word = 8'hC3;
		16'h3C02: out_word = 8'hA0;
		16'h3C03: out_word = 8'h39;
		16'h3C04: out_word = 8'hC3;
		16'h3C05: out_word = 8'h10;
		16'h3C06: out_word = 8'h3C;
		16'h3C07: out_word = 8'hC3;
		16'h3C08: out_word = 8'h10;
		16'h3C09: out_word = 8'h3C;
		16'h3C0A: out_word = 8'hC3;
		16'h3C0B: out_word = 8'h10;
		16'h3C0C: out_word = 8'h3C;
		16'h3C0D: out_word = 8'hC3;
		16'h3C0E: out_word = 8'h10;
		16'h3C0F: out_word = 8'h3C;
		16'h3C10: out_word = 8'h3E;
		16'h3C11: out_word = 8'h7F;
		16'h3C12: out_word = 8'hDB;
		16'h3C13: out_word = 8'hFE;
		16'h3C14: out_word = 8'h1F;
		16'h3C15: out_word = 8'hD8;
		16'h3C16: out_word = 8'h3E;
		16'h3C17: out_word = 8'hFE;
		16'h3C18: out_word = 8'hDB;
		16'h3C19: out_word = 8'hFE;
		16'h3C1A: out_word = 8'h1F;
		16'h3C1B: out_word = 8'hD8;
		16'h3C1C: out_word = 8'h3E;
		16'h3C1D: out_word = 8'h07;
		16'h3C1E: out_word = 8'hD3;
		16'h3C1F: out_word = 8'hFE;
		16'h3C20: out_word = 8'h3E;
		16'h3C21: out_word = 8'h02;
		16'h3C22: out_word = 8'hCD;
		16'h3C23: out_word = 8'h01;
		16'h3C24: out_word = 8'h16;
		16'h3C25: out_word = 8'hAF;
		16'h3C26: out_word = 8'h32;
		16'h3C27: out_word = 8'h3C;
		16'h3C28: out_word = 8'h5C;
		16'h3C29: out_word = 8'h3E;
		16'h3C2A: out_word = 8'h16;
		16'h3C2B: out_word = 8'hD7;
		16'h3C2C: out_word = 8'hAF;
		16'h3C2D: out_word = 8'hD7;
		16'h3C2E: out_word = 8'hAF;
		16'h3C2F: out_word = 8'hD7;
		16'h3C30: out_word = 8'h1E;
		16'h3C31: out_word = 8'h08;
		16'h3C32: out_word = 8'h43;
		16'h3C33: out_word = 8'h50;
		16'h3C34: out_word = 8'h78;
		16'h3C35: out_word = 8'h3D;
		16'h3C36: out_word = 8'hCB;
		16'h3C37: out_word = 8'h17;
		16'h3C38: out_word = 8'hCB;
		16'h3C39: out_word = 8'h17;
		16'h3C3A: out_word = 8'hCB;
		16'h3C3B: out_word = 8'h17;
		16'h3C3C: out_word = 8'h82;
		16'h3C3D: out_word = 8'h3D;
		16'h3C3E: out_word = 8'h32;
		16'h3C3F: out_word = 8'h8F;
		16'h3C40: out_word = 8'h5C;
		16'h3C41: out_word = 8'h21;
		16'h3C42: out_word = 8'h8F;
		16'h3C43: out_word = 8'h3C;
		16'h3C44: out_word = 8'h4B;
		16'h3C45: out_word = 8'h7E;
		16'h3C46: out_word = 8'hD7;
		16'h3C47: out_word = 8'h23;
		16'h3C48: out_word = 8'h0D;
		16'h3C49: out_word = 8'h20;
		16'h3C4A: out_word = 8'hFA;
		16'h3C4B: out_word = 8'h10;
		16'h3C4C: out_word = 8'hE7;
		16'h3C4D: out_word = 8'h43;
		16'h3C4E: out_word = 8'h15;
		16'h3C4F: out_word = 8'h20;
		16'h3C50: out_word = 8'hE3;
		16'h3C51: out_word = 8'h21;
		16'h3C52: out_word = 8'h00;
		16'h3C53: out_word = 8'h48;
		16'h3C54: out_word = 8'h54;
		16'h3C55: out_word = 8'h5D;
		16'h3C56: out_word = 8'h13;
		16'h3C57: out_word = 8'hAF;
		16'h3C58: out_word = 8'h77;
		16'h3C59: out_word = 8'h01;
		16'h3C5A: out_word = 8'hFF;
		16'h3C5B: out_word = 8'h0F;
		16'h3C5C: out_word = 8'hED;
		16'h3C5D: out_word = 8'hB0;
		16'h3C5E: out_word = 8'hEB;
		16'h3C5F: out_word = 8'h11;
		16'h3C60: out_word = 8'h00;
		16'h3C61: out_word = 8'h59;
		16'h3C62: out_word = 8'h01;
		16'h3C63: out_word = 8'h00;
		16'h3C64: out_word = 8'h02;
		16'h3C65: out_word = 8'hED;
		16'h3C66: out_word = 8'hB0;
		16'h3C67: out_word = 8'hF3;
		16'h3C68: out_word = 8'h11;
		16'h3C69: out_word = 8'h70;
		16'h3C6A: out_word = 8'h03;
		16'h3C6B: out_word = 8'h2E;
		16'h3C6C: out_word = 8'h07;
		16'h3C6D: out_word = 8'h01;
		16'h3C6E: out_word = 8'h99;
		16'h3C6F: out_word = 8'h00;
		16'h3C70: out_word = 8'h0B;
		16'h3C71: out_word = 8'h78;
		16'h3C72: out_word = 8'hB1;
		16'h3C73: out_word = 8'h20;
		16'h3C74: out_word = 8'hFB;
		16'h3C75: out_word = 8'h7D;
		16'h3C76: out_word = 8'hEE;
		16'h3C77: out_word = 8'h10;
		16'h3C78: out_word = 8'h6F;
		16'h3C79: out_word = 8'hD3;
		16'h3C7A: out_word = 8'hFE;
		16'h3C7B: out_word = 8'h1B;
		16'h3C7C: out_word = 8'h7A;
		16'h3C7D: out_word = 8'hB3;
		16'h3C7E: out_word = 8'h20;
		16'h3C7F: out_word = 8'hED;
		16'h3C80: out_word = 8'h01;
		16'h3C81: out_word = 8'h00;
		16'h3C82: out_word = 8'h00;
		16'h3C83: out_word = 8'h0B;
		16'h3C84: out_word = 8'h78;
		16'h3C85: out_word = 8'hB1;
		16'h3C86: out_word = 8'h20;
		16'h3C87: out_word = 8'hFB;
		16'h3C88: out_word = 8'h0B;
		16'h3C89: out_word = 8'h78;
		16'h3C8A: out_word = 8'hB1;
		16'h3C8B: out_word = 8'h20;
		16'h3C8C: out_word = 8'hFB;
		16'h3C8D: out_word = 8'h18;
		16'h3C8E: out_word = 8'hD9;
		16'h3C8F: out_word = 8'h13;
		16'h3C90: out_word = 8'h00;
		16'h3C91: out_word = 8'h31;
		16'h3C92: out_word = 8'h39;
		16'h3C93: out_word = 8'h13;
		16'h3C94: out_word = 8'h01;
		16'h3C95: out_word = 8'h38;
		16'h3C96: out_word = 8'h36;
		16'h3C97: out_word = 8'h00;
		16'h3C98: out_word = 8'h00;
		16'h3C99: out_word = 8'h00;
		16'h3C9A: out_word = 8'h00;
		16'h3C9B: out_word = 8'h00;
		16'h3C9C: out_word = 8'h00;
		16'h3C9D: out_word = 8'h00;
		16'h3C9E: out_word = 8'h00;
		16'h3C9F: out_word = 8'h00;
		16'h3CA0: out_word = 8'h00;
		16'h3CA1: out_word = 8'h00;
		16'h3CA2: out_word = 8'h00;
		16'h3CA3: out_word = 8'h00;
		16'h3CA4: out_word = 8'h00;
		16'h3CA5: out_word = 8'h00;
		16'h3CA6: out_word = 8'h00;
		16'h3CA7: out_word = 8'h00;
		16'h3CA8: out_word = 8'h00;
		16'h3CA9: out_word = 8'h00;
		16'h3CAA: out_word = 8'h00;
		16'h3CAB: out_word = 8'h00;
		16'h3CAC: out_word = 8'h00;
		16'h3CAD: out_word = 8'h00;
		16'h3CAE: out_word = 8'h00;
		16'h3CAF: out_word = 8'h00;
		16'h3CB0: out_word = 8'h00;
		16'h3CB1: out_word = 8'h00;
		16'h3CB2: out_word = 8'h00;
		16'h3CB3: out_word = 8'h00;
		16'h3CB4: out_word = 8'h00;
		16'h3CB5: out_word = 8'h00;
		16'h3CB6: out_word = 8'h00;
		16'h3CB7: out_word = 8'h00;
		16'h3CB8: out_word = 8'h00;
		16'h3CB9: out_word = 8'h00;
		16'h3CBA: out_word = 8'h00;
		16'h3CBB: out_word = 8'h00;
		16'h3CBC: out_word = 8'h00;
		16'h3CBD: out_word = 8'h00;
		16'h3CBE: out_word = 8'h00;
		16'h3CBF: out_word = 8'h00;
		16'h3CC0: out_word = 8'h00;
		16'h3CC1: out_word = 8'h00;
		16'h3CC2: out_word = 8'h00;
		16'h3CC3: out_word = 8'h00;
		16'h3CC4: out_word = 8'h00;
		16'h3CC5: out_word = 8'h00;
		16'h3CC6: out_word = 8'h00;
		16'h3CC7: out_word = 8'h00;
		16'h3CC8: out_word = 8'h00;
		16'h3CC9: out_word = 8'h00;
		16'h3CCA: out_word = 8'h00;
		16'h3CCB: out_word = 8'h00;
		16'h3CCC: out_word = 8'h00;
		16'h3CCD: out_word = 8'h00;
		16'h3CCE: out_word = 8'h00;
		16'h3CCF: out_word = 8'h00;
		16'h3CD0: out_word = 8'h00;
		16'h3CD1: out_word = 8'h00;
		16'h3CD2: out_word = 8'h00;
		16'h3CD3: out_word = 8'h00;
		16'h3CD4: out_word = 8'h00;
		16'h3CD5: out_word = 8'h00;
		16'h3CD6: out_word = 8'h00;
		16'h3CD7: out_word = 8'h00;
		16'h3CD8: out_word = 8'h00;
		16'h3CD9: out_word = 8'h00;
		16'h3CDA: out_word = 8'h00;
		16'h3CDB: out_word = 8'h00;
		16'h3CDC: out_word = 8'h00;
		16'h3CDD: out_word = 8'h00;
		16'h3CDE: out_word = 8'h00;
		16'h3CDF: out_word = 8'h00;
		16'h3CE0: out_word = 8'h00;
		16'h3CE1: out_word = 8'h00;
		16'h3CE2: out_word = 8'h00;
		16'h3CE3: out_word = 8'h00;
		16'h3CE4: out_word = 8'h00;
		16'h3CE5: out_word = 8'h00;
		16'h3CE6: out_word = 8'h00;
		16'h3CE7: out_word = 8'h00;
		16'h3CE8: out_word = 8'h00;
		16'h3CE9: out_word = 8'h00;
		16'h3CEA: out_word = 8'h00;
		16'h3CEB: out_word = 8'h00;
		16'h3CEC: out_word = 8'h00;
		16'h3CED: out_word = 8'h00;
		16'h3CEE: out_word = 8'h00;
		16'h3CEF: out_word = 8'h00;
		16'h3CF0: out_word = 8'h00;
		16'h3CF1: out_word = 8'h00;
		16'h3CF2: out_word = 8'h00;
		16'h3CF3: out_word = 8'h00;
		16'h3CF4: out_word = 8'h00;
		16'h3CF5: out_word = 8'h00;
		16'h3CF6: out_word = 8'h00;
		16'h3CF7: out_word = 8'h00;
		16'h3CF8: out_word = 8'h00;
		16'h3CF9: out_word = 8'h00;
		16'h3CFA: out_word = 8'h00;
		16'h3CFB: out_word = 8'h00;
		16'h3CFC: out_word = 8'h00;
		16'h3CFD: out_word = 8'h00;
		16'h3CFE: out_word = 8'h00;
		16'h3CFF: out_word = 8'h00;
		16'h3D00: out_word = 8'h00;
		16'h3D01: out_word = 8'h00;
		16'h3D02: out_word = 8'h00;
		16'h3D03: out_word = 8'h00;
		16'h3D04: out_word = 8'h00;
		16'h3D05: out_word = 8'h00;
		16'h3D06: out_word = 8'h00;
		16'h3D07: out_word = 8'h00;
		16'h3D08: out_word = 8'h00;
		16'h3D09: out_word = 8'h10;
		16'h3D0A: out_word = 8'h10;
		16'h3D0B: out_word = 8'h10;
		16'h3D0C: out_word = 8'h10;
		16'h3D0D: out_word = 8'h00;
		16'h3D0E: out_word = 8'h10;
		16'h3D0F: out_word = 8'h00;
		16'h3D10: out_word = 8'h00;
		16'h3D11: out_word = 8'h24;
		16'h3D12: out_word = 8'h24;
		16'h3D13: out_word = 8'h00;
		16'h3D14: out_word = 8'h00;
		16'h3D15: out_word = 8'h00;
		16'h3D16: out_word = 8'h00;
		16'h3D17: out_word = 8'h00;
		16'h3D18: out_word = 8'h00;
		16'h3D19: out_word = 8'h24;
		16'h3D1A: out_word = 8'h7E;
		16'h3D1B: out_word = 8'h24;
		16'h3D1C: out_word = 8'h24;
		16'h3D1D: out_word = 8'h7E;
		16'h3D1E: out_word = 8'h24;
		16'h3D1F: out_word = 8'h00;
		16'h3D20: out_word = 8'h00;
		16'h3D21: out_word = 8'h08;
		16'h3D22: out_word = 8'h3E;
		16'h3D23: out_word = 8'h28;
		16'h3D24: out_word = 8'h3E;
		16'h3D25: out_word = 8'h0A;
		16'h3D26: out_word = 8'h3E;
		16'h3D27: out_word = 8'h08;
		16'h3D28: out_word = 8'h00;
		16'h3D29: out_word = 8'h62;
		16'h3D2A: out_word = 8'h64;
		16'h3D2B: out_word = 8'h08;
		16'h3D2C: out_word = 8'h10;
		16'h3D2D: out_word = 8'h26;
		16'h3D2E: out_word = 8'h46;
		16'h3D2F: out_word = 8'h00;
		16'h3D30: out_word = 8'h00;
		16'h3D31: out_word = 8'h10;
		16'h3D32: out_word = 8'h28;
		16'h3D33: out_word = 8'h10;
		16'h3D34: out_word = 8'h2A;
		16'h3D35: out_word = 8'h44;
		16'h3D36: out_word = 8'h3A;
		16'h3D37: out_word = 8'h00;
		16'h3D38: out_word = 8'h00;
		16'h3D39: out_word = 8'h08;
		16'h3D3A: out_word = 8'h10;
		16'h3D3B: out_word = 8'h00;
		16'h3D3C: out_word = 8'h00;
		16'h3D3D: out_word = 8'h00;
		16'h3D3E: out_word = 8'h00;
		16'h3D3F: out_word = 8'h00;
		16'h3D40: out_word = 8'h00;
		16'h3D41: out_word = 8'h04;
		16'h3D42: out_word = 8'h08;
		16'h3D43: out_word = 8'h08;
		16'h3D44: out_word = 8'h08;
		16'h3D45: out_word = 8'h08;
		16'h3D46: out_word = 8'h04;
		16'h3D47: out_word = 8'h00;
		16'h3D48: out_word = 8'h00;
		16'h3D49: out_word = 8'h20;
		16'h3D4A: out_word = 8'h10;
		16'h3D4B: out_word = 8'h10;
		16'h3D4C: out_word = 8'h10;
		16'h3D4D: out_word = 8'h10;
		16'h3D4E: out_word = 8'h20;
		16'h3D4F: out_word = 8'h00;
		16'h3D50: out_word = 8'h00;
		16'h3D51: out_word = 8'h00;
		16'h3D52: out_word = 8'h14;
		16'h3D53: out_word = 8'h08;
		16'h3D54: out_word = 8'h3E;
		16'h3D55: out_word = 8'h08;
		16'h3D56: out_word = 8'h14;
		16'h3D57: out_word = 8'h00;
		16'h3D58: out_word = 8'h00;
		16'h3D59: out_word = 8'h00;
		16'h3D5A: out_word = 8'h08;
		16'h3D5B: out_word = 8'h08;
		16'h3D5C: out_word = 8'h3E;
		16'h3D5D: out_word = 8'h08;
		16'h3D5E: out_word = 8'h08;
		16'h3D5F: out_word = 8'h00;
		16'h3D60: out_word = 8'h00;
		16'h3D61: out_word = 8'h00;
		16'h3D62: out_word = 8'h00;
		16'h3D63: out_word = 8'h00;
		16'h3D64: out_word = 8'h00;
		16'h3D65: out_word = 8'h08;
		16'h3D66: out_word = 8'h08;
		16'h3D67: out_word = 8'h10;
		16'h3D68: out_word = 8'h00;
		16'h3D69: out_word = 8'h00;
		16'h3D6A: out_word = 8'h00;
		16'h3D6B: out_word = 8'h00;
		16'h3D6C: out_word = 8'h3E;
		16'h3D6D: out_word = 8'h00;
		16'h3D6E: out_word = 8'h00;
		16'h3D6F: out_word = 8'h00;
		16'h3D70: out_word = 8'h00;
		16'h3D71: out_word = 8'h00;
		16'h3D72: out_word = 8'h00;
		16'h3D73: out_word = 8'h00;
		16'h3D74: out_word = 8'h00;
		16'h3D75: out_word = 8'h18;
		16'h3D76: out_word = 8'h18;
		16'h3D77: out_word = 8'h00;
		16'h3D78: out_word = 8'h00;
		16'h3D79: out_word = 8'h00;
		16'h3D7A: out_word = 8'h02;
		16'h3D7B: out_word = 8'h04;
		16'h3D7C: out_word = 8'h08;
		16'h3D7D: out_word = 8'h10;
		16'h3D7E: out_word = 8'h20;
		16'h3D7F: out_word = 8'h00;
		16'h3D80: out_word = 8'h00;
		16'h3D81: out_word = 8'h3C;
		16'h3D82: out_word = 8'h46;
		16'h3D83: out_word = 8'h4A;
		16'h3D84: out_word = 8'h52;
		16'h3D85: out_word = 8'h62;
		16'h3D86: out_word = 8'h3C;
		16'h3D87: out_word = 8'h00;
		16'h3D88: out_word = 8'h00;
		16'h3D89: out_word = 8'h18;
		16'h3D8A: out_word = 8'h28;
		16'h3D8B: out_word = 8'h08;
		16'h3D8C: out_word = 8'h08;
		16'h3D8D: out_word = 8'h08;
		16'h3D8E: out_word = 8'h3E;
		16'h3D8F: out_word = 8'h00;
		16'h3D90: out_word = 8'h00;
		16'h3D91: out_word = 8'h3C;
		16'h3D92: out_word = 8'h42;
		16'h3D93: out_word = 8'h02;
		16'h3D94: out_word = 8'h3C;
		16'h3D95: out_word = 8'h40;
		16'h3D96: out_word = 8'h7E;
		16'h3D97: out_word = 8'h00;
		16'h3D98: out_word = 8'h00;
		16'h3D99: out_word = 8'h3C;
		16'h3D9A: out_word = 8'h42;
		16'h3D9B: out_word = 8'h0C;
		16'h3D9C: out_word = 8'h02;
		16'h3D9D: out_word = 8'h42;
		16'h3D9E: out_word = 8'h3C;
		16'h3D9F: out_word = 8'h00;
		16'h3DA0: out_word = 8'h00;
		16'h3DA1: out_word = 8'h08;
		16'h3DA2: out_word = 8'h18;
		16'h3DA3: out_word = 8'h28;
		16'h3DA4: out_word = 8'h48;
		16'h3DA5: out_word = 8'h7E;
		16'h3DA6: out_word = 8'h08;
		16'h3DA7: out_word = 8'h00;
		16'h3DA8: out_word = 8'h00;
		16'h3DA9: out_word = 8'h7E;
		16'h3DAA: out_word = 8'h40;
		16'h3DAB: out_word = 8'h7C;
		16'h3DAC: out_word = 8'h02;
		16'h3DAD: out_word = 8'h42;
		16'h3DAE: out_word = 8'h3C;
		16'h3DAF: out_word = 8'h00;
		16'h3DB0: out_word = 8'h00;
		16'h3DB1: out_word = 8'h3C;
		16'h3DB2: out_word = 8'h40;
		16'h3DB3: out_word = 8'h7C;
		16'h3DB4: out_word = 8'h42;
		16'h3DB5: out_word = 8'h42;
		16'h3DB6: out_word = 8'h3C;
		16'h3DB7: out_word = 8'h00;
		16'h3DB8: out_word = 8'h00;
		16'h3DB9: out_word = 8'h7E;
		16'h3DBA: out_word = 8'h02;
		16'h3DBB: out_word = 8'h04;
		16'h3DBC: out_word = 8'h08;
		16'h3DBD: out_word = 8'h10;
		16'h3DBE: out_word = 8'h10;
		16'h3DBF: out_word = 8'h00;
		16'h3DC0: out_word = 8'h00;
		16'h3DC1: out_word = 8'h3C;
		16'h3DC2: out_word = 8'h42;
		16'h3DC3: out_word = 8'h3C;
		16'h3DC4: out_word = 8'h42;
		16'h3DC5: out_word = 8'h42;
		16'h3DC6: out_word = 8'h3C;
		16'h3DC7: out_word = 8'h00;
		16'h3DC8: out_word = 8'h00;
		16'h3DC9: out_word = 8'h3C;
		16'h3DCA: out_word = 8'h42;
		16'h3DCB: out_word = 8'h42;
		16'h3DCC: out_word = 8'h3E;
		16'h3DCD: out_word = 8'h02;
		16'h3DCE: out_word = 8'h3C;
		16'h3DCF: out_word = 8'h00;
		16'h3DD0: out_word = 8'h00;
		16'h3DD1: out_word = 8'h00;
		16'h3DD2: out_word = 8'h00;
		16'h3DD3: out_word = 8'h10;
		16'h3DD4: out_word = 8'h00;
		16'h3DD5: out_word = 8'h00;
		16'h3DD6: out_word = 8'h10;
		16'h3DD7: out_word = 8'h00;
		16'h3DD8: out_word = 8'h00;
		16'h3DD9: out_word = 8'h00;
		16'h3DDA: out_word = 8'h10;
		16'h3DDB: out_word = 8'h00;
		16'h3DDC: out_word = 8'h00;
		16'h3DDD: out_word = 8'h10;
		16'h3DDE: out_word = 8'h10;
		16'h3DDF: out_word = 8'h20;
		16'h3DE0: out_word = 8'h00;
		16'h3DE1: out_word = 8'h00;
		16'h3DE2: out_word = 8'h04;
		16'h3DE3: out_word = 8'h08;
		16'h3DE4: out_word = 8'h10;
		16'h3DE5: out_word = 8'h08;
		16'h3DE6: out_word = 8'h04;
		16'h3DE7: out_word = 8'h00;
		16'h3DE8: out_word = 8'h00;
		16'h3DE9: out_word = 8'h00;
		16'h3DEA: out_word = 8'h00;
		16'h3DEB: out_word = 8'h3E;
		16'h3DEC: out_word = 8'h00;
		16'h3DED: out_word = 8'h3E;
		16'h3DEE: out_word = 8'h00;
		16'h3DEF: out_word = 8'h00;
		16'h3DF0: out_word = 8'h00;
		16'h3DF1: out_word = 8'h00;
		16'h3DF2: out_word = 8'h10;
		16'h3DF3: out_word = 8'h08;
		16'h3DF4: out_word = 8'h04;
		16'h3DF5: out_word = 8'h08;
		16'h3DF6: out_word = 8'h10;
		16'h3DF7: out_word = 8'h00;
		16'h3DF8: out_word = 8'h00;
		16'h3DF9: out_word = 8'h3C;
		16'h3DFA: out_word = 8'h42;
		16'h3DFB: out_word = 8'h04;
		16'h3DFC: out_word = 8'h08;
		16'h3DFD: out_word = 8'h00;
		16'h3DFE: out_word = 8'h08;
		16'h3DFF: out_word = 8'h00;
		16'h3E00: out_word = 8'h00;
		16'h3E01: out_word = 8'h3C;
		16'h3E02: out_word = 8'h4A;
		16'h3E03: out_word = 8'h56;
		16'h3E04: out_word = 8'h5E;
		16'h3E05: out_word = 8'h40;
		16'h3E06: out_word = 8'h3C;
		16'h3E07: out_word = 8'h00;
		16'h3E08: out_word = 8'h00;
		16'h3E09: out_word = 8'h3C;
		16'h3E0A: out_word = 8'h42;
		16'h3E0B: out_word = 8'h42;
		16'h3E0C: out_word = 8'h7E;
		16'h3E0D: out_word = 8'h42;
		16'h3E0E: out_word = 8'h42;
		16'h3E0F: out_word = 8'h00;
		16'h3E10: out_word = 8'h00;
		16'h3E11: out_word = 8'h7C;
		16'h3E12: out_word = 8'h42;
		16'h3E13: out_word = 8'h7C;
		16'h3E14: out_word = 8'h42;
		16'h3E15: out_word = 8'h42;
		16'h3E16: out_word = 8'h7C;
		16'h3E17: out_word = 8'h00;
		16'h3E18: out_word = 8'h00;
		16'h3E19: out_word = 8'h3C;
		16'h3E1A: out_word = 8'h42;
		16'h3E1B: out_word = 8'h40;
		16'h3E1C: out_word = 8'h40;
		16'h3E1D: out_word = 8'h42;
		16'h3E1E: out_word = 8'h3C;
		16'h3E1F: out_word = 8'h00;
		16'h3E20: out_word = 8'h00;
		16'h3E21: out_word = 8'h78;
		16'h3E22: out_word = 8'h44;
		16'h3E23: out_word = 8'h42;
		16'h3E24: out_word = 8'h42;
		16'h3E25: out_word = 8'h44;
		16'h3E26: out_word = 8'h78;
		16'h3E27: out_word = 8'h00;
		16'h3E28: out_word = 8'h00;
		16'h3E29: out_word = 8'h7E;
		16'h3E2A: out_word = 8'h40;
		16'h3E2B: out_word = 8'h7C;
		16'h3E2C: out_word = 8'h40;
		16'h3E2D: out_word = 8'h40;
		16'h3E2E: out_word = 8'h7E;
		16'h3E2F: out_word = 8'h00;
		16'h3E30: out_word = 8'h00;
		16'h3E31: out_word = 8'h7E;
		16'h3E32: out_word = 8'h40;
		16'h3E33: out_word = 8'h7C;
		16'h3E34: out_word = 8'h40;
		16'h3E35: out_word = 8'h40;
		16'h3E36: out_word = 8'h40;
		16'h3E37: out_word = 8'h00;
		16'h3E38: out_word = 8'h00;
		16'h3E39: out_word = 8'h3C;
		16'h3E3A: out_word = 8'h42;
		16'h3E3B: out_word = 8'h40;
		16'h3E3C: out_word = 8'h4E;
		16'h3E3D: out_word = 8'h42;
		16'h3E3E: out_word = 8'h3C;
		16'h3E3F: out_word = 8'h00;
		16'h3E40: out_word = 8'h00;
		16'h3E41: out_word = 8'h42;
		16'h3E42: out_word = 8'h42;
		16'h3E43: out_word = 8'h7E;
		16'h3E44: out_word = 8'h42;
		16'h3E45: out_word = 8'h42;
		16'h3E46: out_word = 8'h42;
		16'h3E47: out_word = 8'h00;
		16'h3E48: out_word = 8'h00;
		16'h3E49: out_word = 8'h3E;
		16'h3E4A: out_word = 8'h08;
		16'h3E4B: out_word = 8'h08;
		16'h3E4C: out_word = 8'h08;
		16'h3E4D: out_word = 8'h08;
		16'h3E4E: out_word = 8'h3E;
		16'h3E4F: out_word = 8'h00;
		16'h3E50: out_word = 8'h00;
		16'h3E51: out_word = 8'h02;
		16'h3E52: out_word = 8'h02;
		16'h3E53: out_word = 8'h02;
		16'h3E54: out_word = 8'h42;
		16'h3E55: out_word = 8'h42;
		16'h3E56: out_word = 8'h3C;
		16'h3E57: out_word = 8'h00;
		16'h3E58: out_word = 8'h00;
		16'h3E59: out_word = 8'h44;
		16'h3E5A: out_word = 8'h48;
		16'h3E5B: out_word = 8'h70;
		16'h3E5C: out_word = 8'h48;
		16'h3E5D: out_word = 8'h44;
		16'h3E5E: out_word = 8'h42;
		16'h3E5F: out_word = 8'h00;
		16'h3E60: out_word = 8'h00;
		16'h3E61: out_word = 8'h40;
		16'h3E62: out_word = 8'h40;
		16'h3E63: out_word = 8'h40;
		16'h3E64: out_word = 8'h40;
		16'h3E65: out_word = 8'h40;
		16'h3E66: out_word = 8'h7E;
		16'h3E67: out_word = 8'h00;
		16'h3E68: out_word = 8'h00;
		16'h3E69: out_word = 8'h42;
		16'h3E6A: out_word = 8'h66;
		16'h3E6B: out_word = 8'h5A;
		16'h3E6C: out_word = 8'h42;
		16'h3E6D: out_word = 8'h42;
		16'h3E6E: out_word = 8'h42;
		16'h3E6F: out_word = 8'h00;
		16'h3E70: out_word = 8'h00;
		16'h3E71: out_word = 8'h42;
		16'h3E72: out_word = 8'h62;
		16'h3E73: out_word = 8'h52;
		16'h3E74: out_word = 8'h4A;
		16'h3E75: out_word = 8'h46;
		16'h3E76: out_word = 8'h42;
		16'h3E77: out_word = 8'h00;
		16'h3E78: out_word = 8'h00;
		16'h3E79: out_word = 8'h3C;
		16'h3E7A: out_word = 8'h42;
		16'h3E7B: out_word = 8'h42;
		16'h3E7C: out_word = 8'h42;
		16'h3E7D: out_word = 8'h42;
		16'h3E7E: out_word = 8'h3C;
		16'h3E7F: out_word = 8'h00;
		16'h3E80: out_word = 8'h00;
		16'h3E81: out_word = 8'h7C;
		16'h3E82: out_word = 8'h42;
		16'h3E83: out_word = 8'h42;
		16'h3E84: out_word = 8'h7C;
		16'h3E85: out_word = 8'h40;
		16'h3E86: out_word = 8'h40;
		16'h3E87: out_word = 8'h00;
		16'h3E88: out_word = 8'h00;
		16'h3E89: out_word = 8'h3C;
		16'h3E8A: out_word = 8'h42;
		16'h3E8B: out_word = 8'h42;
		16'h3E8C: out_word = 8'h52;
		16'h3E8D: out_word = 8'h4A;
		16'h3E8E: out_word = 8'h3C;
		16'h3E8F: out_word = 8'h00;
		16'h3E90: out_word = 8'h00;
		16'h3E91: out_word = 8'h7C;
		16'h3E92: out_word = 8'h42;
		16'h3E93: out_word = 8'h42;
		16'h3E94: out_word = 8'h7C;
		16'h3E95: out_word = 8'h44;
		16'h3E96: out_word = 8'h42;
		16'h3E97: out_word = 8'h00;
		16'h3E98: out_word = 8'h00;
		16'h3E99: out_word = 8'h3C;
		16'h3E9A: out_word = 8'h40;
		16'h3E9B: out_word = 8'h3C;
		16'h3E9C: out_word = 8'h02;
		16'h3E9D: out_word = 8'h42;
		16'h3E9E: out_word = 8'h3C;
		16'h3E9F: out_word = 8'h00;
		16'h3EA0: out_word = 8'h00;
		16'h3EA1: out_word = 8'hFE;
		16'h3EA2: out_word = 8'h10;
		16'h3EA3: out_word = 8'h10;
		16'h3EA4: out_word = 8'h10;
		16'h3EA5: out_word = 8'h10;
		16'h3EA6: out_word = 8'h10;
		16'h3EA7: out_word = 8'h00;
		16'h3EA8: out_word = 8'h00;
		16'h3EA9: out_word = 8'h42;
		16'h3EAA: out_word = 8'h42;
		16'h3EAB: out_word = 8'h42;
		16'h3EAC: out_word = 8'h42;
		16'h3EAD: out_word = 8'h42;
		16'h3EAE: out_word = 8'h3C;
		16'h3EAF: out_word = 8'h00;
		16'h3EB0: out_word = 8'h00;
		16'h3EB1: out_word = 8'h42;
		16'h3EB2: out_word = 8'h42;
		16'h3EB3: out_word = 8'h42;
		16'h3EB4: out_word = 8'h42;
		16'h3EB5: out_word = 8'h24;
		16'h3EB6: out_word = 8'h18;
		16'h3EB7: out_word = 8'h00;
		16'h3EB8: out_word = 8'h00;
		16'h3EB9: out_word = 8'h42;
		16'h3EBA: out_word = 8'h42;
		16'h3EBB: out_word = 8'h42;
		16'h3EBC: out_word = 8'h42;
		16'h3EBD: out_word = 8'h5A;
		16'h3EBE: out_word = 8'h24;
		16'h3EBF: out_word = 8'h00;
		16'h3EC0: out_word = 8'h00;
		16'h3EC1: out_word = 8'h42;
		16'h3EC2: out_word = 8'h24;
		16'h3EC3: out_word = 8'h18;
		16'h3EC4: out_word = 8'h18;
		16'h3EC5: out_word = 8'h24;
		16'h3EC6: out_word = 8'h42;
		16'h3EC7: out_word = 8'h00;
		16'h3EC8: out_word = 8'h00;
		16'h3EC9: out_word = 8'h82;
		16'h3ECA: out_word = 8'h44;
		16'h3ECB: out_word = 8'h28;
		16'h3ECC: out_word = 8'h10;
		16'h3ECD: out_word = 8'h10;
		16'h3ECE: out_word = 8'h10;
		16'h3ECF: out_word = 8'h00;
		16'h3ED0: out_word = 8'h00;
		16'h3ED1: out_word = 8'h7E;
		16'h3ED2: out_word = 8'h04;
		16'h3ED3: out_word = 8'h08;
		16'h3ED4: out_word = 8'h10;
		16'h3ED5: out_word = 8'h20;
		16'h3ED6: out_word = 8'h7E;
		16'h3ED7: out_word = 8'h00;
		16'h3ED8: out_word = 8'h00;
		16'h3ED9: out_word = 8'h0E;
		16'h3EDA: out_word = 8'h08;
		16'h3EDB: out_word = 8'h08;
		16'h3EDC: out_word = 8'h08;
		16'h3EDD: out_word = 8'h08;
		16'h3EDE: out_word = 8'h0E;
		16'h3EDF: out_word = 8'h00;
		16'h3EE0: out_word = 8'h00;
		16'h3EE1: out_word = 8'h00;
		16'h3EE2: out_word = 8'h40;
		16'h3EE3: out_word = 8'h20;
		16'h3EE4: out_word = 8'h10;
		16'h3EE5: out_word = 8'h08;
		16'h3EE6: out_word = 8'h04;
		16'h3EE7: out_word = 8'h00;
		16'h3EE8: out_word = 8'h00;
		16'h3EE9: out_word = 8'h70;
		16'h3EEA: out_word = 8'h10;
		16'h3EEB: out_word = 8'h10;
		16'h3EEC: out_word = 8'h10;
		16'h3EED: out_word = 8'h10;
		16'h3EEE: out_word = 8'h70;
		16'h3EEF: out_word = 8'h00;
		16'h3EF0: out_word = 8'h00;
		16'h3EF1: out_word = 8'h10;
		16'h3EF2: out_word = 8'h38;
		16'h3EF3: out_word = 8'h54;
		16'h3EF4: out_word = 8'h10;
		16'h3EF5: out_word = 8'h10;
		16'h3EF6: out_word = 8'h10;
		16'h3EF7: out_word = 8'h00;
		16'h3EF8: out_word = 8'h00;
		16'h3EF9: out_word = 8'h00;
		16'h3EFA: out_word = 8'h00;
		16'h3EFB: out_word = 8'h00;
		16'h3EFC: out_word = 8'h00;
		16'h3EFD: out_word = 8'h00;
		16'h3EFE: out_word = 8'h00;
		16'h3EFF: out_word = 8'hFF;
		16'h3F00: out_word = 8'h00;
		16'h3F01: out_word = 8'h1C;
		16'h3F02: out_word = 8'h22;
		16'h3F03: out_word = 8'h78;
		16'h3F04: out_word = 8'h20;
		16'h3F05: out_word = 8'h20;
		16'h3F06: out_word = 8'h7E;
		16'h3F07: out_word = 8'h00;
		16'h3F08: out_word = 8'h00;
		16'h3F09: out_word = 8'h00;
		16'h3F0A: out_word = 8'h38;
		16'h3F0B: out_word = 8'h04;
		16'h3F0C: out_word = 8'h3C;
		16'h3F0D: out_word = 8'h44;
		16'h3F0E: out_word = 8'h3C;
		16'h3F0F: out_word = 8'h00;
		16'h3F10: out_word = 8'h00;
		16'h3F11: out_word = 8'h20;
		16'h3F12: out_word = 8'h20;
		16'h3F13: out_word = 8'h3C;
		16'h3F14: out_word = 8'h22;
		16'h3F15: out_word = 8'h22;
		16'h3F16: out_word = 8'h3C;
		16'h3F17: out_word = 8'h00;
		16'h3F18: out_word = 8'h00;
		16'h3F19: out_word = 8'h00;
		16'h3F1A: out_word = 8'h1C;
		16'h3F1B: out_word = 8'h20;
		16'h3F1C: out_word = 8'h20;
		16'h3F1D: out_word = 8'h20;
		16'h3F1E: out_word = 8'h1C;
		16'h3F1F: out_word = 8'h00;
		16'h3F20: out_word = 8'h00;
		16'h3F21: out_word = 8'h04;
		16'h3F22: out_word = 8'h04;
		16'h3F23: out_word = 8'h3C;
		16'h3F24: out_word = 8'h44;
		16'h3F25: out_word = 8'h44;
		16'h3F26: out_word = 8'h3C;
		16'h3F27: out_word = 8'h00;
		16'h3F28: out_word = 8'h00;
		16'h3F29: out_word = 8'h00;
		16'h3F2A: out_word = 8'h38;
		16'h3F2B: out_word = 8'h44;
		16'h3F2C: out_word = 8'h78;
		16'h3F2D: out_word = 8'h40;
		16'h3F2E: out_word = 8'h3C;
		16'h3F2F: out_word = 8'h00;
		16'h3F30: out_word = 8'h00;
		16'h3F31: out_word = 8'h0C;
		16'h3F32: out_word = 8'h10;
		16'h3F33: out_word = 8'h18;
		16'h3F34: out_word = 8'h10;
		16'h3F35: out_word = 8'h10;
		16'h3F36: out_word = 8'h10;
		16'h3F37: out_word = 8'h00;
		16'h3F38: out_word = 8'h00;
		16'h3F39: out_word = 8'h00;
		16'h3F3A: out_word = 8'h3C;
		16'h3F3B: out_word = 8'h44;
		16'h3F3C: out_word = 8'h44;
		16'h3F3D: out_word = 8'h3C;
		16'h3F3E: out_word = 8'h04;
		16'h3F3F: out_word = 8'h38;
		16'h3F40: out_word = 8'h00;
		16'h3F41: out_word = 8'h40;
		16'h3F42: out_word = 8'h40;
		16'h3F43: out_word = 8'h78;
		16'h3F44: out_word = 8'h44;
		16'h3F45: out_word = 8'h44;
		16'h3F46: out_word = 8'h44;
		16'h3F47: out_word = 8'h00;
		16'h3F48: out_word = 8'h00;
		16'h3F49: out_word = 8'h10;
		16'h3F4A: out_word = 8'h00;
		16'h3F4B: out_word = 8'h30;
		16'h3F4C: out_word = 8'h10;
		16'h3F4D: out_word = 8'h10;
		16'h3F4E: out_word = 8'h38;
		16'h3F4F: out_word = 8'h00;
		16'h3F50: out_word = 8'h00;
		16'h3F51: out_word = 8'h04;
		16'h3F52: out_word = 8'h00;
		16'h3F53: out_word = 8'h04;
		16'h3F54: out_word = 8'h04;
		16'h3F55: out_word = 8'h04;
		16'h3F56: out_word = 8'h24;
		16'h3F57: out_word = 8'h18;
		16'h3F58: out_word = 8'h00;
		16'h3F59: out_word = 8'h20;
		16'h3F5A: out_word = 8'h28;
		16'h3F5B: out_word = 8'h30;
		16'h3F5C: out_word = 8'h30;
		16'h3F5D: out_word = 8'h28;
		16'h3F5E: out_word = 8'h24;
		16'h3F5F: out_word = 8'h00;
		16'h3F60: out_word = 8'h00;
		16'h3F61: out_word = 8'h10;
		16'h3F62: out_word = 8'h10;
		16'h3F63: out_word = 8'h10;
		16'h3F64: out_word = 8'h10;
		16'h3F65: out_word = 8'h10;
		16'h3F66: out_word = 8'h0C;
		16'h3F67: out_word = 8'h00;
		16'h3F68: out_word = 8'h00;
		16'h3F69: out_word = 8'h00;
		16'h3F6A: out_word = 8'h68;
		16'h3F6B: out_word = 8'h54;
		16'h3F6C: out_word = 8'h54;
		16'h3F6D: out_word = 8'h54;
		16'h3F6E: out_word = 8'h54;
		16'h3F6F: out_word = 8'h00;
		16'h3F70: out_word = 8'h00;
		16'h3F71: out_word = 8'h00;
		16'h3F72: out_word = 8'h78;
		16'h3F73: out_word = 8'h44;
		16'h3F74: out_word = 8'h44;
		16'h3F75: out_word = 8'h44;
		16'h3F76: out_word = 8'h44;
		16'h3F77: out_word = 8'h00;
		16'h3F78: out_word = 8'h00;
		16'h3F79: out_word = 8'h00;
		16'h3F7A: out_word = 8'h38;
		16'h3F7B: out_word = 8'h44;
		16'h3F7C: out_word = 8'h44;
		16'h3F7D: out_word = 8'h44;
		16'h3F7E: out_word = 8'h38;
		16'h3F7F: out_word = 8'h00;
		16'h3F80: out_word = 8'h00;
		16'h3F81: out_word = 8'h00;
		16'h3F82: out_word = 8'h78;
		16'h3F83: out_word = 8'h44;
		16'h3F84: out_word = 8'h44;
		16'h3F85: out_word = 8'h78;
		16'h3F86: out_word = 8'h40;
		16'h3F87: out_word = 8'h40;
		16'h3F88: out_word = 8'h00;
		16'h3F89: out_word = 8'h00;
		16'h3F8A: out_word = 8'h3C;
		16'h3F8B: out_word = 8'h44;
		16'h3F8C: out_word = 8'h44;
		16'h3F8D: out_word = 8'h3C;
		16'h3F8E: out_word = 8'h04;
		16'h3F8F: out_word = 8'h06;
		16'h3F90: out_word = 8'h00;
		16'h3F91: out_word = 8'h00;
		16'h3F92: out_word = 8'h1C;
		16'h3F93: out_word = 8'h20;
		16'h3F94: out_word = 8'h20;
		16'h3F95: out_word = 8'h20;
		16'h3F96: out_word = 8'h20;
		16'h3F97: out_word = 8'h00;
		16'h3F98: out_word = 8'h00;
		16'h3F99: out_word = 8'h00;
		16'h3F9A: out_word = 8'h38;
		16'h3F9B: out_word = 8'h40;
		16'h3F9C: out_word = 8'h38;
		16'h3F9D: out_word = 8'h04;
		16'h3F9E: out_word = 8'h78;
		16'h3F9F: out_word = 8'h00;
		16'h3FA0: out_word = 8'h00;
		16'h3FA1: out_word = 8'h10;
		16'h3FA2: out_word = 8'h38;
		16'h3FA3: out_word = 8'h10;
		16'h3FA4: out_word = 8'h10;
		16'h3FA5: out_word = 8'h10;
		16'h3FA6: out_word = 8'h0C;
		16'h3FA7: out_word = 8'h00;
		16'h3FA8: out_word = 8'h00;
		16'h3FA9: out_word = 8'h00;
		16'h3FAA: out_word = 8'h44;
		16'h3FAB: out_word = 8'h44;
		16'h3FAC: out_word = 8'h44;
		16'h3FAD: out_word = 8'h44;
		16'h3FAE: out_word = 8'h38;
		16'h3FAF: out_word = 8'h00;
		16'h3FB0: out_word = 8'h00;
		16'h3FB1: out_word = 8'h00;
		16'h3FB2: out_word = 8'h44;
		16'h3FB3: out_word = 8'h44;
		16'h3FB4: out_word = 8'h28;
		16'h3FB5: out_word = 8'h28;
		16'h3FB6: out_word = 8'h10;
		16'h3FB7: out_word = 8'h00;
		16'h3FB8: out_word = 8'h00;
		16'h3FB9: out_word = 8'h00;
		16'h3FBA: out_word = 8'h44;
		16'h3FBB: out_word = 8'h54;
		16'h3FBC: out_word = 8'h54;
		16'h3FBD: out_word = 8'h54;
		16'h3FBE: out_word = 8'h28;
		16'h3FBF: out_word = 8'h00;
		16'h3FC0: out_word = 8'h00;
		16'h3FC1: out_word = 8'h00;
		16'h3FC2: out_word = 8'h44;
		16'h3FC3: out_word = 8'h28;
		16'h3FC4: out_word = 8'h10;
		16'h3FC5: out_word = 8'h28;
		16'h3FC6: out_word = 8'h44;
		16'h3FC7: out_word = 8'h00;
		16'h3FC8: out_word = 8'h00;
		16'h3FC9: out_word = 8'h00;
		16'h3FCA: out_word = 8'h44;
		16'h3FCB: out_word = 8'h44;
		16'h3FCC: out_word = 8'h44;
		16'h3FCD: out_word = 8'h3C;
		16'h3FCE: out_word = 8'h04;
		16'h3FCF: out_word = 8'h38;
		16'h3FD0: out_word = 8'h00;
		16'h3FD1: out_word = 8'h00;
		16'h3FD2: out_word = 8'h7C;
		16'h3FD3: out_word = 8'h08;
		16'h3FD4: out_word = 8'h10;
		16'h3FD5: out_word = 8'h20;
		16'h3FD6: out_word = 8'h7C;
		16'h3FD7: out_word = 8'h00;
		16'h3FD8: out_word = 8'h00;
		16'h3FD9: out_word = 8'h0E;
		16'h3FDA: out_word = 8'h08;
		16'h3FDB: out_word = 8'h30;
		16'h3FDC: out_word = 8'h08;
		16'h3FDD: out_word = 8'h08;
		16'h3FDE: out_word = 8'h0E;
		16'h3FDF: out_word = 8'h00;
		16'h3FE0: out_word = 8'h00;
		16'h3FE1: out_word = 8'h08;
		16'h3FE2: out_word = 8'h08;
		16'h3FE3: out_word = 8'h08;
		16'h3FE4: out_word = 8'h08;
		16'h3FE5: out_word = 8'h08;
		16'h3FE6: out_word = 8'h08;
		16'h3FE7: out_word = 8'h00;
		16'h3FE8: out_word = 8'h00;
		16'h3FE9: out_word = 8'h70;
		16'h3FEA: out_word = 8'h10;
		16'h3FEB: out_word = 8'h0C;
		16'h3FEC: out_word = 8'h10;
		16'h3FED: out_word = 8'h10;
		16'h3FEE: out_word = 8'h70;
		16'h3FEF: out_word = 8'h00;
		16'h3FF0: out_word = 8'h00;
		16'h3FF1: out_word = 8'h14;
		16'h3FF2: out_word = 8'h28;
		16'h3FF3: out_word = 8'h00;
		16'h3FF4: out_word = 8'h00;
		16'h3FF5: out_word = 8'h00;
		16'h3FF6: out_word = 8'h00;
		16'h3FF7: out_word = 8'h00;
		16'h3FF8: out_word = 8'h3C;
		16'h3FF9: out_word = 8'h42;
		16'h3FFA: out_word = 8'h99;
		16'h3FFB: out_word = 8'hA1;
		16'h3FFC: out_word = 8'hA1;
		16'h3FFD: out_word = 8'h99;
		16'h3FFE: out_word = 8'h42;
		16'h3FFF: out_word = 8'h3C;
		16'h4000: out_word = 8'hF3;
		16'h4001: out_word = 8'h11;
		16'h4002: out_word = 8'hFF;
		16'h4003: out_word = 8'hFF;
		16'h4004: out_word = 8'hC3;
		16'h4005: out_word = 8'h50;
		16'h4006: out_word = 8'h3C;
		16'h4007: out_word = 8'h01;
		16'h4008: out_word = 8'h00;
		16'h4009: out_word = 8'hD3;
		16'h400A: out_word = 8'hFE;
		16'h400B: out_word = 8'h3E;
		16'h400C: out_word = 8'h3F;
		16'h400D: out_word = 8'h18;
		16'h400E: out_word = 8'h04;
		16'h400F: out_word = 8'h00;
		16'h4010: out_word = 8'hC3;
		16'h4011: out_word = 8'h82;
		16'h4012: out_word = 8'h3D;
		16'h4013: out_word = 8'hED;
		16'h4014: out_word = 8'h47;
		16'h4015: out_word = 8'hC3;
		16'h4016: out_word = 8'h1B;
		16'h4017: out_word = 8'h00;
		16'h4018: out_word = 8'hC3;
		16'h4019: out_word = 8'h07;
		16'h401A: out_word = 8'h27;
		16'h401B: out_word = 8'h00;
		16'h401C: out_word = 8'h00;
		16'h401D: out_word = 8'h00;
		16'h401E: out_word = 8'h18;
		16'h401F: out_word = 8'h04;
		16'h4020: out_word = 8'hC3;
		16'h4021: out_word = 8'h72;
		16'h4022: out_word = 8'h2F;
		16'h4023: out_word = 8'hC9;
		16'h4024: out_word = 8'h62;
		16'h4025: out_word = 8'h6B;
		16'h4026: out_word = 8'h18;
		16'h4027: out_word = 8'h03;
		16'h4028: out_word = 8'hC3;
		16'h4029: out_word = 8'h23;
		16'h402A: out_word = 8'h23;
		16'h402B: out_word = 8'hAF;
		16'h402C: out_word = 8'h47;
		16'h402D: out_word = 8'h4F;
		16'h402E: out_word = 8'hF9;
		16'h402F: out_word = 8'h18;
		16'h4030: out_word = 8'h09;
		16'h4031: out_word = 8'hFF;
		16'h4032: out_word = 8'hFF;
		16'h4033: out_word = 8'hFF;
		16'h4034: out_word = 8'hFF;
		16'h4035: out_word = 8'hFF;
		16'h4036: out_word = 8'hFF;
		16'h4037: out_word = 8'hFF;
		16'h4038: out_word = 8'hFB;
		16'h4039: out_word = 8'hC9;
		16'h403A: out_word = 8'hC5;
		16'h403B: out_word = 8'hC5;
		16'h403C: out_word = 8'hC5;
		16'h403D: out_word = 8'hC5;
		16'h403E: out_word = 8'hC5;
		16'h403F: out_word = 8'hC5;
		16'h4040: out_word = 8'hC5;
		16'h4041: out_word = 8'hC5;
		16'h4042: out_word = 8'h21;
		16'h4043: out_word = 8'h00;
		16'h4044: out_word = 8'hA5;
		16'h4045: out_word = 8'h39;
		16'h4046: out_word = 8'h38;
		16'h4047: out_word = 8'hF2;
		16'h4048: out_word = 8'h22;
		16'h4049: out_word = 8'hB4;
		16'h404A: out_word = 8'h5C;
		16'h404B: out_word = 8'h11;
		16'h404C: out_word = 8'hAF;
		16'h404D: out_word = 8'h3E;
		16'h404E: out_word = 8'h01;
		16'h404F: out_word = 8'hA8;
		16'h4050: out_word = 8'h00;
		16'h4051: out_word = 8'h7B;
		16'h4052: out_word = 8'hEB;
		16'h4053: out_word = 8'h31;
		16'h4054: out_word = 8'h00;
		16'h4055: out_word = 8'h60;
		16'h4056: out_word = 8'h22;
		16'h4057: out_word = 8'h00;
		16'h4058: out_word = 8'h5F;
		16'h4059: out_word = 8'h21;
		16'h405A: out_word = 8'h79;
		16'h405B: out_word = 8'h00;
		16'h405C: out_word = 8'hE5;
		16'h405D: out_word = 8'h21;
		16'h405E: out_word = 8'h2F;
		16'h405F: out_word = 8'h3D;
		16'h4060: out_word = 8'hE5;
		16'h4061: out_word = 8'h21;
		16'h4062: out_word = 8'hED;
		16'h4063: out_word = 8'hB8;
		16'h4064: out_word = 8'h18;
		16'h4065: out_word = 8'h03;
		16'h4066: out_word = 8'hC3;
		16'h4067: out_word = 8'h56;
		16'h4068: out_word = 8'h2A;
		16'h4069: out_word = 8'h22;
		16'h406A: out_word = 8'h10;
		16'h406B: out_word = 8'h5F;
		16'h406C: out_word = 8'hF5;
		16'h406D: out_word = 8'h3E;
		16'h406E: out_word = 8'hC9;
		16'h406F: out_word = 8'h32;
		16'h4070: out_word = 8'h12;
		16'h4071: out_word = 8'h5F;
		16'h4072: out_word = 8'hF1;
		16'h4073: out_word = 8'h2A;
		16'h4074: out_word = 8'h00;
		16'h4075: out_word = 8'h5F;
		16'h4076: out_word = 8'hC3;
		16'h4077: out_word = 8'h10;
		16'h4078: out_word = 8'h5F;
		16'h4079: out_word = 8'hEB;
		16'h407A: out_word = 8'h23;
		16'h407B: out_word = 8'h22;
		16'h407C: out_word = 8'h7B;
		16'h407D: out_word = 8'h5C;
		16'h407E: out_word = 8'h2B;
		16'h407F: out_word = 8'h01;
		16'h4080: out_word = 8'h40;
		16'h4081: out_word = 8'h05;
		16'h4082: out_word = 8'hED;
		16'h4083: out_word = 8'h43;
		16'h4084: out_word = 8'h38;
		16'h4085: out_word = 8'h5C;
		16'h4086: out_word = 8'h22;
		16'h4087: out_word = 8'hB2;
		16'h4088: out_word = 8'h5C;
		16'h4089: out_word = 8'h21;
		16'h408A: out_word = 8'h00;
		16'h408B: out_word = 8'h3C;
		16'h408C: out_word = 8'h22;
		16'h408D: out_word = 8'h36;
		16'h408E: out_word = 8'h5C;
		16'h408F: out_word = 8'h2A;
		16'h4090: out_word = 8'hB2;
		16'h4091: out_word = 8'h5C;
		16'h4092: out_word = 8'h36;
		16'h4093: out_word = 8'h3E;
		16'h4094: out_word = 8'h2B;
		16'h4095: out_word = 8'hF9;
		16'h4096: out_word = 8'h2B;
		16'h4097: out_word = 8'h2B;
		16'h4098: out_word = 8'h22;
		16'h4099: out_word = 8'h3D;
		16'h409A: out_word = 8'h5C;
		16'h409B: out_word = 8'h11;
		16'h409C: out_word = 8'h03;
		16'h409D: out_word = 8'h13;
		16'h409E: out_word = 8'hD5;
		16'h409F: out_word = 8'hED;
		16'h40A0: out_word = 8'h56;
		16'h40A1: out_word = 8'hFD;
		16'h40A2: out_word = 8'h21;
		16'h40A3: out_word = 8'h3A;
		16'h40A4: out_word = 8'h5C;
		16'h40A5: out_word = 8'h21;
		16'h40A6: out_word = 8'hB6;
		16'h40A7: out_word = 8'h5C;
		16'h40A8: out_word = 8'h22;
		16'h40A9: out_word = 8'h4F;
		16'h40AA: out_word = 8'h5C;
		16'h40AB: out_word = 8'h11;
		16'h40AC: out_word = 8'hAF;
		16'h40AD: out_word = 8'h15;
		16'h40AE: out_word = 8'h01;
		16'h40AF: out_word = 8'h15;
		16'h40B0: out_word = 8'h00;
		16'h40B1: out_word = 8'hEB;
		16'h40B2: out_word = 8'hCD;
		16'h40B3: out_word = 8'h17;
		16'h40B4: out_word = 8'h01;
		16'h40B5: out_word = 8'hEB;
		16'h40B6: out_word = 8'h2B;
		16'h40B7: out_word = 8'h22;
		16'h40B8: out_word = 8'h57;
		16'h40B9: out_word = 8'h5C;
		16'h40BA: out_word = 8'h23;
		16'h40BB: out_word = 8'h22;
		16'h40BC: out_word = 8'h53;
		16'h40BD: out_word = 8'h5C;
		16'h40BE: out_word = 8'h22;
		16'h40BF: out_word = 8'h4B;
		16'h40C0: out_word = 8'h5C;
		16'h40C1: out_word = 8'h36;
		16'h40C2: out_word = 8'h80;
		16'h40C3: out_word = 8'h23;
		16'h40C4: out_word = 8'h22;
		16'h40C5: out_word = 8'h59;
		16'h40C6: out_word = 8'h5C;
		16'h40C7: out_word = 8'h36;
		16'h40C8: out_word = 8'h0D;
		16'h40C9: out_word = 8'h23;
		16'h40CA: out_word = 8'h36;
		16'h40CB: out_word = 8'h80;
		16'h40CC: out_word = 8'h23;
		16'h40CD: out_word = 8'h22;
		16'h40CE: out_word = 8'h61;
		16'h40CF: out_word = 8'h5C;
		16'h40D0: out_word = 8'h22;
		16'h40D1: out_word = 8'h63;
		16'h40D2: out_word = 8'h5C;
		16'h40D3: out_word = 8'h22;
		16'h40D4: out_word = 8'h65;
		16'h40D5: out_word = 8'h5C;
		16'h40D6: out_word = 8'h3E;
		16'h40D7: out_word = 8'h38;
		16'h40D8: out_word = 8'h32;
		16'h40D9: out_word = 8'h8D;
		16'h40DA: out_word = 8'h5C;
		16'h40DB: out_word = 8'h32;
		16'h40DC: out_word = 8'h8F;
		16'h40DD: out_word = 8'h5C;
		16'h40DE: out_word = 8'h32;
		16'h40DF: out_word = 8'h48;
		16'h40E0: out_word = 8'h5C;
		16'h40E1: out_word = 8'h21;
		16'h40E2: out_word = 8'h23;
		16'h40E3: out_word = 8'h02;
		16'h40E4: out_word = 8'h22;
		16'h40E5: out_word = 8'h09;
		16'h40E6: out_word = 8'h5C;
		16'h40E7: out_word = 8'hFD;
		16'h40E8: out_word = 8'h35;
		16'h40E9: out_word = 8'hC6;
		16'h40EA: out_word = 8'hFD;
		16'h40EB: out_word = 8'h35;
		16'h40EC: out_word = 8'hCA;
		16'h40ED: out_word = 8'h21;
		16'h40EE: out_word = 8'hC6;
		16'h40EF: out_word = 8'h15;
		16'h40F0: out_word = 8'h11;
		16'h40F1: out_word = 8'h10;
		16'h40F2: out_word = 8'h5C;
		16'h40F3: out_word = 8'h01;
		16'h40F4: out_word = 8'h0E;
		16'h40F5: out_word = 8'h00;
		16'h40F6: out_word = 8'hCD;
		16'h40F7: out_word = 8'h17;
		16'h40F8: out_word = 8'h01;
		16'h40F9: out_word = 8'hFD;
		16'h40FA: out_word = 8'hCB;
		16'h40FB: out_word = 8'h01;
		16'h40FC: out_word = 8'hCE;
		16'h40FD: out_word = 8'h21;
		16'h40FE: out_word = 8'hC2;
		16'h40FF: out_word = 8'h5C;
		16'h4100: out_word = 8'h36;
		16'h4101: out_word = 8'hC9;
		16'h4102: out_word = 8'hE7;
		16'h4103: out_word = 8'hDF;
		16'h4104: out_word = 8'h0E;
		16'h4105: out_word = 8'h21;
		16'h4106: out_word = 8'h6B;
		16'h4107: out_word = 8'h5C;
		16'h4108: out_word = 8'h36;
		16'h4109: out_word = 8'h02;
		16'h410A: out_word = 8'h21;
		16'h410B: out_word = 8'h8B;
		16'h410C: out_word = 8'h12;
		16'h410D: out_word = 8'hE5;
		16'h410E: out_word = 8'h3E;
		16'h410F: out_word = 8'hAA;
		16'h4110: out_word = 8'h32;
		16'h4111: out_word = 8'h81;
		16'h4112: out_word = 8'h5C;
		16'h4113: out_word = 8'hFB;
		16'h4114: out_word = 8'hC3;
		16'h4115: out_word = 8'h31;
		16'h4116: out_word = 8'h3D;
		16'h4117: out_word = 8'h22;
		16'h4118: out_word = 8'h00;
		16'h4119: out_word = 8'h5F;
		16'h411A: out_word = 8'h21;
		16'h411B: out_word = 8'h2F;
		16'h411C: out_word = 8'h3D;
		16'h411D: out_word = 8'hE5;
		16'h411E: out_word = 8'h21;
		16'h411F: out_word = 8'hED;
		16'h4120: out_word = 8'hB0;
		16'h4121: out_word = 8'h22;
		16'h4122: out_word = 8'h10;
		16'h4123: out_word = 8'h5F;
		16'h4124: out_word = 8'h2A;
		16'h4125: out_word = 8'h00;
		16'h4126: out_word = 8'h5F;
		16'h4127: out_word = 8'hC3;
		16'h4128: out_word = 8'h10;
		16'h4129: out_word = 8'h5F;
		16'h412A: out_word = 8'hCD;
		16'h412B: out_word = 8'hE5;
		16'h412C: out_word = 8'h20;
		16'h412D: out_word = 8'hCD;
		16'h412E: out_word = 8'h97;
		16'h412F: out_word = 8'h1D;
		16'h4130: out_word = 8'h2A;
		16'h4131: out_word = 8'h59;
		16'h4132: out_word = 8'h5C;
		16'h4133: out_word = 8'h23;
		16'h4134: out_word = 8'h5E;
		16'h4135: out_word = 8'h23;
		16'h4136: out_word = 8'h56;
		16'h4137: out_word = 8'h7A;
		16'h4138: out_word = 8'hB3;
		16'h4139: out_word = 8'hEB;
		16'h413A: out_word = 8'h28;
		16'h413B: out_word = 8'h04;
		16'h413C: out_word = 8'hAF;
		16'h413D: out_word = 8'h32;
		16'h413E: out_word = 8'h10;
		16'h413F: out_word = 8'h5D;
		16'h4140: out_word = 8'hE5;
		16'h4141: out_word = 8'hCD;
		16'h4142: out_word = 8'h32;
		16'h4143: out_word = 8'h02;
		16'h4144: out_word = 8'hE1;
		16'h4145: out_word = 8'h22;
		16'h4146: out_word = 8'h42;
		16'h4147: out_word = 8'h5C;
		16'h4148: out_word = 8'hAF;
		16'h4149: out_word = 8'h32;
		16'h414A: out_word = 8'h44;
		16'h414B: out_word = 8'h5C;
		16'h414C: out_word = 8'hE7;
		16'h414D: out_word = 8'hB0;
		16'h414E: out_word = 8'h16;
		16'h414F: out_word = 8'h2A;
		16'h4150: out_word = 8'h53;
		16'h4151: out_word = 8'h5C;
		16'h4152: out_word = 8'h2B;
		16'h4153: out_word = 8'h22;
		16'h4154: out_word = 8'h57;
		16'h4155: out_word = 8'h5C;
		16'h4156: out_word = 8'hED;
		16'h4157: out_word = 8'h7B;
		16'h4158: out_word = 8'h3D;
		16'h4159: out_word = 8'h5C;
		16'h415A: out_word = 8'h3A;
		16'h415B: out_word = 8'h10;
		16'h415C: out_word = 8'h5D;
		16'h415D: out_word = 8'hB7;
		16'h415E: out_word = 8'h21;
		16'h415F: out_word = 8'h76;
		16'h4160: out_word = 8'h1B;
		16'h4161: out_word = 8'h28;
		16'h4162: out_word = 8'h03;
		16'h4163: out_word = 8'hE7;
		16'h4164: out_word = 8'hB0;
		16'h4165: out_word = 8'h1B;
		16'h4166: out_word = 8'hE5;
		16'h4167: out_word = 8'h21;
		16'h4168: out_word = 8'hC2;
		16'h4169: out_word = 8'h5C;
		16'h416A: out_word = 8'hE5;
		16'h416B: out_word = 8'hC9;
		16'h416C: out_word = 8'hCD;
		16'h416D: out_word = 8'hF1;
		16'h416E: out_word = 8'h20;
		16'h416F: out_word = 8'hCD;
		16'h4170: out_word = 8'h4A;
		16'h4171: out_word = 8'h29;
		16'h4172: out_word = 8'h3E;
		16'h4173: out_word = 8'hFF;
		16'h4174: out_word = 8'h32;
		16'h4175: out_word = 8'h15;
		16'h4176: out_word = 8'h5D;
		16'h4177: out_word = 8'hAF;
		16'h4178: out_word = 8'h32;
		16'h4179: out_word = 8'hF7;
		16'h417A: out_word = 8'h5C;
		16'h417B: out_word = 8'h3E;
		16'h417C: out_word = 8'hAA;
		16'h417D: out_word = 8'h32;
		16'h417E: out_word = 8'h17;
		16'h417F: out_word = 8'h5D;
		16'h4180: out_word = 8'h21;
		16'h4181: out_word = 8'h01;
		16'h4182: out_word = 8'h02;
		16'h4183: out_word = 8'h22;
		16'h4184: out_word = 8'h1A;
		16'h4185: out_word = 8'h5D;
		16'h4186: out_word = 8'h21;
		16'h4187: out_word = 8'h00;
		16'h4188: out_word = 8'h00;
		16'h4189: out_word = 8'h39;
		16'h418A: out_word = 8'h22;
		16'h418B: out_word = 8'h1C;
		16'h418C: out_word = 8'h5D;
		16'h418D: out_word = 8'h2B;
		16'h418E: out_word = 8'h2B;
		16'h418F: out_word = 8'hF9;
		16'h4190: out_word = 8'hCD;
		16'h4191: out_word = 8'h1D;
		16'h4192: out_word = 8'h02;
		16'h4193: out_word = 8'h2A;
		16'h4194: out_word = 8'hB2;
		16'h4195: out_word = 8'h5C;
		16'h4196: out_word = 8'hED;
		16'h4197: out_word = 8'h5B;
		16'h4198: out_word = 8'h5D;
		16'h4199: out_word = 8'h5C;
		16'h419A: out_word = 8'hED;
		16'h419B: out_word = 8'h52;
		16'h419C: out_word = 8'hEB;
		16'h419D: out_word = 8'h30;
		16'h419E: out_word = 8'h06;
		16'h419F: out_word = 8'hB7;
		16'h41A0: out_word = 8'h11;
		16'h41A1: out_word = 8'h01;
		16'h41A2: out_word = 8'h01;
		16'h41A3: out_word = 8'hED;
		16'h41A4: out_word = 8'h52;
		16'h41A5: out_word = 8'h22;
		16'h41A6: out_word = 8'h5D;
		16'h41A7: out_word = 8'h5C;
		16'h41A8: out_word = 8'hCD;
		16'h41A9: out_word = 8'hC7;
		16'h41AA: out_word = 8'h01;
		16'h41AB: out_word = 8'hCA;
		16'h41AC: out_word = 8'hD3;
		16'h41AD: out_word = 8'h01;
		16'h41AE: out_word = 8'hFE;
		16'h41AF: out_word = 8'hEA;
		16'h41B0: out_word = 8'h23;
		16'h41B1: out_word = 8'h20;
		16'h41B2: out_word = 8'hF5;
		16'h41B3: out_word = 8'hCD;
		16'h41B4: out_word = 8'hC7;
		16'h41B5: out_word = 8'h01;
		16'h41B6: out_word = 8'h28;
		16'h41B7: out_word = 8'hF3;
		16'h41B8: out_word = 8'hFE;
		16'h41B9: out_word = 8'h3A;
		16'h41BA: out_word = 8'hC2;
		16'h41BB: out_word = 8'hD3;
		16'h41BC: out_word = 8'h01;
		16'h41BD: out_word = 8'h23;
		16'h41BE: out_word = 8'hCD;
		16'h41BF: out_word = 8'h48;
		16'h41C0: out_word = 8'h30;
		16'h41C1: out_word = 8'h2A;
		16'h41C2: out_word = 8'h11;
		16'h41C3: out_word = 8'h5D;
		16'h41C4: out_word = 8'hC3;
		16'h41C5: out_word = 8'h0A;
		16'h41C6: out_word = 8'h03;
		16'h41C7: out_word = 8'h7E;
		16'h41C8: out_word = 8'hFE;
		16'h41C9: out_word = 8'h0D;
		16'h41CA: out_word = 8'hC8;
		16'h41CB: out_word = 8'hFE;
		16'h41CC: out_word = 8'h80;
		16'h41CD: out_word = 8'hC8;
		16'h41CE: out_word = 8'hB7;
		16'h41CF: out_word = 8'hC9;
		16'h41D0: out_word = 8'hCD;
		16'h41D1: out_word = 8'h43;
		16'h41D2: out_word = 8'h1E;
		16'h41D3: out_word = 8'h21;
		16'h41D4: out_word = 8'h00;
		16'h41D5: out_word = 8'h00;
		16'h41D6: out_word = 8'h22;
		16'h41D7: out_word = 8'hF8;
		16'h41D8: out_word = 8'h5C;
		16'h41D9: out_word = 8'hCD;
		16'h41DA: out_word = 8'hE5;
		16'h41DB: out_word = 8'h20;
		16'h41DC: out_word = 8'hCD;
		16'h41DD: out_word = 8'h63;
		16'h41DE: out_word = 8'h1D;
		16'h41DF: out_word = 8'h21;
		16'h41E0: out_word = 8'h17;
		16'h41E1: out_word = 8'h5D;
		16'h41E2: out_word = 8'h36;
		16'h41E3: out_word = 8'hAA;
		16'h41E4: out_word = 8'h21;
		16'h41E5: out_word = 8'h1F;
		16'h41E6: out_word = 8'h5D;
		16'h41E7: out_word = 8'h7E;
		16'h41E8: out_word = 8'hB7;
		16'h41E9: out_word = 8'h36;
		16'h41EA: out_word = 8'h00;
		16'h41EB: out_word = 8'h20;
		16'h41EC: out_word = 8'h06;
		16'h41ED: out_word = 8'hCD;
		16'h41EE: out_word = 8'h1C;
		16'h41EF: out_word = 8'h1E;
		16'h41F0: out_word = 8'hCD;
		16'h41F1: out_word = 8'h12;
		16'h41F2: out_word = 8'h02;
		16'h41F3: out_word = 8'hED;
		16'h41F4: out_word = 8'h7B;
		16'h41F5: out_word = 8'h1C;
		16'h41F6: out_word = 8'h5D;
		16'h41F7: out_word = 8'h2A;
		16'h41F8: out_word = 8'h1A;
		16'h41F9: out_word = 8'h5D;
		16'h41FA: out_word = 8'hED;
		16'h41FB: out_word = 8'h4B;
		16'h41FC: out_word = 8'h0F;
		16'h41FD: out_word = 8'h5D;
		16'h41FE: out_word = 8'h06;
		16'h41FF: out_word = 8'h00;
		16'h4200: out_word = 8'hE9;
		16'h4201: out_word = 8'hCD;
		16'h4202: out_word = 8'h32;
		16'h4203: out_word = 8'h02;
		16'h4204: out_word = 8'hFD;
		16'h4205: out_word = 8'hCB;
		16'h4206: out_word = 8'h00;
		16'h4207: out_word = 8'h7E;
		16'h4208: out_word = 8'hC0;
		16'h4209: out_word = 8'h11;
		16'h420A: out_word = 8'hC2;
		16'h420B: out_word = 8'h5C;
		16'h420C: out_word = 8'hED;
		16'h420D: out_word = 8'h7B;
		16'h420E: out_word = 8'h3D;
		16'h420F: out_word = 8'h5C;
		16'h4210: out_word = 8'hD5;
		16'h4211: out_word = 8'hC9;
		16'h4212: out_word = 8'hCD;
		16'h4213: out_word = 8'h8C;
		16'h4214: out_word = 8'h1D;
		16'h4215: out_word = 8'hFE;
		16'h4216: out_word = 8'h0D;
		16'h4217: out_word = 8'hC8;
		16'h4218: out_word = 8'hCD;
		16'h4219: out_word = 8'h2A;
		16'h421A: out_word = 8'h1E;
		16'h421B: out_word = 8'h18;
		16'h421C: out_word = 8'hF5;
		16'h421D: out_word = 8'h2A;
		16'h421E: out_word = 8'h3D;
		16'h421F: out_word = 8'h5C;
		16'h4220: out_word = 8'h22;
		16'h4221: out_word = 8'h13;
		16'h4222: out_word = 8'h5D;
		16'h4223: out_word = 8'h2A;
		16'h4224: out_word = 8'h1C;
		16'h4225: out_word = 8'h5D;
		16'h4226: out_word = 8'h2B;
		16'h4227: out_word = 8'h2B;
		16'h4228: out_word = 8'h22;
		16'h4229: out_word = 8'h3D;
		16'h422A: out_word = 8'h5C;
		16'h422B: out_word = 8'h11;
		16'h422C: out_word = 8'h16;
		16'h422D: out_word = 8'h3D;
		16'h422E: out_word = 8'h73;
		16'h422F: out_word = 8'h23;
		16'h4230: out_word = 8'h72;
		16'h4231: out_word = 8'hC9;
		16'h4232: out_word = 8'h2A;
		16'h4233: out_word = 8'h13;
		16'h4234: out_word = 8'h5D;
		16'h4235: out_word = 8'h22;
		16'h4236: out_word = 8'h3D;
		16'h4237: out_word = 8'h5C;
		16'h4238: out_word = 8'hC9;
		16'h4239: out_word = 8'h21;
		16'h423A: out_word = 8'h00;
		16'h423B: out_word = 8'h00;
		16'h423C: out_word = 8'h22;
		16'h423D: out_word = 8'hF7;
		16'h423E: out_word = 8'h5C;
		16'h423F: out_word = 8'h39;
		16'h4240: out_word = 8'h22;
		16'h4241: out_word = 8'h1C;
		16'h4242: out_word = 8'h5D;
		16'h4243: out_word = 8'h2B;
		16'h4244: out_word = 8'h2B;
		16'h4245: out_word = 8'hF9;
		16'h4246: out_word = 8'hCD;
		16'h4247: out_word = 8'h1C;
		16'h4248: out_word = 8'h32;
		16'h4249: out_word = 8'h21;
		16'h424A: out_word = 8'h17;
		16'h424B: out_word = 8'h5D;
		16'h424C: out_word = 8'h7E;
		16'h424D: out_word = 8'hFE;
		16'h424E: out_word = 8'hAA;
		16'h424F: out_word = 8'h3E;
		16'h4250: out_word = 8'h00;
		16'h4251: out_word = 8'h32;
		16'h4252: out_word = 8'h0F;
		16'h4253: out_word = 8'h5D;
		16'h4254: out_word = 8'hCA;
		16'h4255: out_word = 8'hCB;
		16'h4256: out_word = 8'h02;
		16'h4257: out_word = 8'h36;
		16'h4258: out_word = 8'hAA;
		16'h4259: out_word = 8'hCD;
		16'h425A: out_word = 8'h97;
		16'h425B: out_word = 8'h1D;
		16'h425C: out_word = 8'hCD;
		16'h425D: out_word = 8'h88;
		16'h425E: out_word = 8'h1D;
		16'h425F: out_word = 8'h21;
		16'h4260: out_word = 8'h60;
		16'h4261: out_word = 8'h03;
		16'h4262: out_word = 8'hDF;
		16'h4263: out_word = 8'hCD;
		16'h4264: out_word = 8'h9C;
		16'h4265: out_word = 8'h39;
		16'h4266: out_word = 8'h00;
		16'h4267: out_word = 8'hCD;
		16'h4268: out_word = 8'h37;
		16'h4269: out_word = 8'h38;
		16'h426A: out_word = 8'hFB;
		16'h426B: out_word = 8'h20;
		16'h426C: out_word = 8'h04;
		16'h426D: out_word = 8'h21;
		16'h426E: out_word = 8'h00;
		16'h426F: out_word = 8'h10;
		16'h4270: out_word = 8'hDF;
		16'h4271: out_word = 8'h3A;
		16'h4272: out_word = 8'h81;
		16'h4273: out_word = 8'h5C;
		16'h4274: out_word = 8'hFE;
		16'h4275: out_word = 8'hAA;
		16'h4276: out_word = 8'h20;
		16'h4277: out_word = 8'h53;
		16'h4278: out_word = 8'hCD;
		16'h4279: out_word = 8'hF1;
		16'h427A: out_word = 8'h20;
		16'h427B: out_word = 8'h2A;
		16'h427C: out_word = 8'h59;
		16'h427D: out_word = 8'h5C;
		16'h427E: out_word = 8'h3E;
		16'h427F: out_word = 8'hFE;
		16'h4280: out_word = 8'h32;
		16'h4281: out_word = 8'h0E;
		16'h4282: out_word = 8'h5D;
		16'h4283: out_word = 8'h36;
		16'h4284: out_word = 8'hF7;
		16'h4285: out_word = 8'h23;
		16'h4286: out_word = 8'h36;
		16'h4287: out_word = 8'h22;
		16'h4288: out_word = 8'h23;
		16'h4289: out_word = 8'h36;
		16'h428A: out_word = 8'h62;
		16'h428B: out_word = 8'h23;
		16'h428C: out_word = 8'h36;
		16'h428D: out_word = 8'h6F;
		16'h428E: out_word = 8'h23;
		16'h428F: out_word = 8'h36;
		16'h4290: out_word = 8'h6F;
		16'h4291: out_word = 8'h23;
		16'h4292: out_word = 8'h36;
		16'h4293: out_word = 8'h74;
		16'h4294: out_word = 8'h23;
		16'h4295: out_word = 8'h36;
		16'h4296: out_word = 8'h22;
		16'h4297: out_word = 8'h23;
		16'h4298: out_word = 8'h22;
		16'h4299: out_word = 8'h5B;
		16'h429A: out_word = 8'h5C;
		16'h429B: out_word = 8'h36;
		16'h429C: out_word = 8'h0D;
		16'h429D: out_word = 8'h23;
		16'h429E: out_word = 8'h36;
		16'h429F: out_word = 8'h80;
		16'h42A0: out_word = 8'h23;
		16'h42A1: out_word = 8'h22;
		16'h42A2: out_word = 8'h61;
		16'h42A3: out_word = 8'h5C;
		16'h42A4: out_word = 8'h22;
		16'h42A5: out_word = 8'h63;
		16'h42A6: out_word = 8'h5C;
		16'h42A7: out_word = 8'h22;
		16'h42A8: out_word = 8'h65;
		16'h42A9: out_word = 8'h5C;
		16'h42AA: out_word = 8'hFD;
		16'h42AB: out_word = 8'hCB;
		16'h42AC: out_word = 8'h01;
		16'h42AD: out_word = 8'hDE;
		16'h42AE: out_word = 8'h18;
		16'h42AF: out_word = 8'h3F;
		16'h42B0: out_word = 8'h06;
		16'h42B1: out_word = 8'h03;
		16'h42B2: out_word = 8'h7E;
		16'h42B3: out_word = 8'h12;
		16'h42B4: out_word = 8'h23;
		16'h42B5: out_word = 8'h13;
		16'h42B6: out_word = 8'h10;
		16'h42B7: out_word = 8'hFA;
		16'h42B8: out_word = 8'hC9;
		16'h42B9: out_word = 8'h06;
		16'h42BA: out_word = 8'h20;
		16'h42BB: out_word = 8'hC5;
		16'h42BC: out_word = 8'hEE;
		16'h42BD: out_word = 8'h08;
		16'h42BE: out_word = 8'hD3;
		16'h42BF: out_word = 8'hFF;
		16'h42C0: out_word = 8'hF5;
		16'h42C1: out_word = 8'h3E;
		16'h42C2: out_word = 8'h05;
		16'h42C3: out_word = 8'hCD;
		16'h42C4: out_word = 8'hFF;
		16'h42C5: out_word = 8'h3D;
		16'h42C6: out_word = 8'hF1;
		16'h42C7: out_word = 8'hC1;
		16'h42C8: out_word = 8'h10;
		16'h42C9: out_word = 8'hF1;
		16'h42CA: out_word = 8'hC9;
		16'h42CB: out_word = 8'h2A;
		16'h42CC: out_word = 8'h1C;
		16'h42CD: out_word = 8'h5D;
		16'h42CE: out_word = 8'h2B;
		16'h42CF: out_word = 8'h2B;
		16'h42D0: out_word = 8'hF9;
		16'h42D1: out_word = 8'hCD;
		16'h42D2: out_word = 8'hF1;
		16'h42D3: out_word = 8'h20;
		16'h42D4: out_word = 8'hCD;
		16'h42D5: out_word = 8'h83;
		16'h42D6: out_word = 8'h1D;
		16'h42D7: out_word = 8'h3A;
		16'h42D8: out_word = 8'h16;
		16'h42D9: out_word = 8'h5D;
		16'h42DA: out_word = 8'hF6;
		16'h42DB: out_word = 8'h03;
		16'h42DC: out_word = 8'hCD;
		16'h42DD: out_word = 8'hB9;
		16'h42DE: out_word = 8'h02;
		16'h42DF: out_word = 8'h3A;
		16'h42E0: out_word = 8'h16;
		16'h42E1: out_word = 8'h5D;
		16'h42E2: out_word = 8'hCD;
		16'h42E3: out_word = 8'hB9;
		16'h42E4: out_word = 8'h02;
		16'h42E5: out_word = 8'hAF;
		16'h42E6: out_word = 8'h32;
		16'h42E7: out_word = 8'h15;
		16'h42E8: out_word = 8'h5D;
		16'h42E9: out_word = 8'hCD;
		16'h42EA: out_word = 8'h35;
		16'h42EB: out_word = 8'h21;
		16'h42EC: out_word = 8'hCD;
		16'h42ED: out_word = 8'h32;
		16'h42EE: out_word = 8'h30;
		16'h42EF: out_word = 8'hCD;
		16'h42F0: out_word = 8'h9F;
		16'h42F1: out_word = 8'h1D;
		16'h42F2: out_word = 8'h21;
		16'h42F3: out_word = 8'hCB;
		16'h42F4: out_word = 8'h02;
		16'h42F5: out_word = 8'h22;
		16'h42F6: out_word = 8'h1A;
		16'h42F7: out_word = 8'h5D;
		16'h42F8: out_word = 8'hAF;
		16'h42F9: out_word = 8'h32;
		16'h42FA: out_word = 8'h0F;
		16'h42FB: out_word = 8'h5D;
		16'h42FC: out_word = 8'h2A;
		16'h42FD: out_word = 8'h59;
		16'h42FE: out_word = 8'h5C;
		16'h42FF: out_word = 8'hE5;
		16'h4300: out_word = 8'h11;
		16'h4301: out_word = 8'h20;
		16'h4302: out_word = 8'h5D;
		16'h4303: out_word = 8'hCD;
		16'h4304: out_word = 8'hB0;
		16'h4305: out_word = 8'h02;
		16'h4306: out_word = 8'hE1;
		16'h4307: out_word = 8'h22;
		16'h4308: out_word = 8'h11;
		16'h4309: out_word = 8'h5D;
		16'h430A: out_word = 8'h7E;
		16'h430B: out_word = 8'h47;
		16'h430C: out_word = 8'hE6;
		16'h430D: out_word = 8'h80;
		16'h430E: out_word = 8'h78;
		16'h430F: out_word = 8'h28;
		16'h4310: out_word = 8'h09;
		16'h4311: out_word = 8'hFE;
		16'h4312: out_word = 8'hFE;
		16'h4313: out_word = 8'h28;
		16'h4314: out_word = 8'h05;
		16'h4315: out_word = 8'hF5;
		16'h4316: out_word = 8'hCD;
		16'h4317: out_word = 8'hC8;
		16'h4318: out_word = 8'h3D;
		16'h4319: out_word = 8'hF1;
		16'h431A: out_word = 8'h21;
		16'h431B: out_word = 8'hF3;
		16'h431C: out_word = 8'h2F;
		16'h431D: out_word = 8'h2B;
		16'h431E: out_word = 8'h0E;
		16'h431F: out_word = 8'h00;
		16'h4320: out_word = 8'h0C;
		16'h4321: out_word = 8'h57;
		16'h4322: out_word = 8'h3E;
		16'h4323: out_word = 8'h15;
		16'h4324: out_word = 8'hB9;
		16'h4325: out_word = 8'hDA;
		16'h4326: out_word = 8'hD3;
		16'h4327: out_word = 8'h01;
		16'h4328: out_word = 8'h7A;
		16'h4329: out_word = 8'h23;
		16'h432A: out_word = 8'hBE;
		16'h432B: out_word = 8'h20;
		16'h432C: out_word = 8'hF3;
		16'h432D: out_word = 8'hFE;
		16'h432E: out_word = 8'hFE;
		16'h432F: out_word = 8'hC4;
		16'h4330: out_word = 8'h4A;
		16'h4331: out_word = 8'h29;
		16'h4332: out_word = 8'h3E;
		16'h4333: out_word = 8'h09;
		16'h4334: out_word = 8'h32;
		16'h4335: out_word = 8'h06;
		16'h4336: out_word = 8'h5D;
		16'h4337: out_word = 8'hAF;
		16'h4338: out_word = 8'h32;
		16'h4339: out_word = 8'h0F;
		16'h433A: out_word = 8'h5D;
		16'h433B: out_word = 8'h32;
		16'h433C: out_word = 8'hD6;
		16'h433D: out_word = 8'h5C;
		16'h433E: out_word = 8'h32;
		16'h433F: out_word = 8'h10;
		16'h4340: out_word = 8'h5D;
		16'h4341: out_word = 8'h21;
		16'h4342: out_word = 8'h3B;
		16'h4343: out_word = 8'h5C;
		16'h4344: out_word = 8'hCB;
		16'h4345: out_word = 8'hBE;
		16'h4346: out_word = 8'h06;
		16'h4347: out_word = 8'h00;
		16'h4348: out_word = 8'h21;
		16'h4349: out_word = 8'h08;
		16'h434A: out_word = 8'h30;
		16'h434B: out_word = 8'h0D;
		16'h434C: out_word = 8'hCB;
		16'h434D: out_word = 8'h21;
		16'h434E: out_word = 8'h09;
		16'h434F: out_word = 8'h5E;
		16'h4350: out_word = 8'h23;
		16'h4351: out_word = 8'h56;
		16'h4352: out_word = 8'hEB;
		16'h4353: out_word = 8'hE5;
		16'h4354: out_word = 8'h11;
		16'h4355: out_word = 8'h59;
		16'h4356: out_word = 8'h03;
		16'h4357: out_word = 8'hD5;
		16'h4358: out_word = 8'hE9;
		16'h4359: out_word = 8'h21;
		16'h435A: out_word = 8'h3B;
		16'h435B: out_word = 8'h5C;
		16'h435C: out_word = 8'hCB;
		16'h435D: out_word = 8'hFE;
		16'h435E: out_word = 8'hE1;
		16'h435F: out_word = 8'hE9;
		16'h4360: out_word = 8'h16;
		16'h4361: out_word = 8'h01;
		16'h4362: out_word = 8'h05;
		16'h4363: out_word = 8'h2A;
		16'h4364: out_word = 8'h20;
		16'h4365: out_word = 8'h54;
		16'h4366: out_word = 8'h52;
		16'h4367: out_word = 8'h2D;
		16'h4368: out_word = 8'h44;
		16'h4369: out_word = 8'h4F;
		16'h436A: out_word = 8'h53;
		16'h436B: out_word = 8'h20;
		16'h436C: out_word = 8'h56;
		16'h436D: out_word = 8'h65;
		16'h436E: out_word = 8'h72;
		16'h436F: out_word = 8'h20;
		16'h4370: out_word = 8'h36;
		16'h4371: out_word = 8'h2E;
		16'h4372: out_word = 8'h31;
		16'h4373: out_word = 8'h32;
		16'h4374: out_word = 8'h45;
		16'h4375: out_word = 8'h2A;
		16'h4376: out_word = 8'h0D;
		16'h4377: out_word = 8'h0D;
		16'h4378: out_word = 8'h31;
		16'h4379: out_word = 8'h39;
		16'h437A: out_word = 8'h39;
		16'h437B: out_word = 8'h39;
		16'h437C: out_word = 8'h20;
		16'h437D: out_word = 8'h43;
		16'h437E: out_word = 8'h6F;
		16'h437F: out_word = 8'h6D;
		16'h4380: out_word = 8'h70;
		16'h4381: out_word = 8'h6F;
		16'h4382: out_word = 8'h57;
		16'h4383: out_word = 8'h65;
		16'h4384: out_word = 8'h6C;
		16'h4385: out_word = 8'h6C;
		16'h4386: out_word = 8'h63;
		16'h4387: out_word = 8'h6F;
		16'h4388: out_word = 8'h6D;
		16'h4389: out_word = 8'h65;
		16'h438A: out_word = 8'h2C;
		16'h438B: out_word = 8'h20;
		16'h438C: out_word = 8'h32;
		16'h438D: out_word = 8'h30;
		16'h438E: out_word = 8'h30;
		16'h438F: out_word = 8'h35;
		16'h4390: out_word = 8'h20;
		16'h4391: out_word = 8'h41;
		16'h4392: out_word = 8'h6C;
		16'h4393: out_word = 8'h6F;
		16'h4394: out_word = 8'h6E;
		16'h4395: out_word = 8'h65;
		16'h4396: out_word = 8'h2E;
		16'h4397: out_word = 8'h16;
		16'h4398: out_word = 8'h05;
		16'h4399: out_word = 8'h0B;
		16'h439A: out_word = 8'h52;
		16'h439B: out_word = 8'h79;
		16'h439C: out_word = 8'h61;
		16'h439D: out_word = 8'h7A;
		16'h439E: out_word = 8'h61;
		16'h439F: out_word = 8'h6E;
		16'h43A0: out_word = 8'h16;
		16'h43A1: out_word = 8'h07;
		16'h43A2: out_word = 8'h05;
		16'h43A3: out_word = 8'h42;
		16'h43A4: out_word = 8'h45;
		16'h43A5: out_word = 8'h54;
		16'h43A6: out_word = 8'h41;
		16'h43A7: out_word = 8'h31;
		16'h43A8: out_word = 8'h30;
		16'h43A9: out_word = 8'h32;
		16'h43AA: out_word = 8'h34;
		16'h43AB: out_word = 8'h00;
		16'h43AC: out_word = 8'hCD;
		16'h43AD: out_word = 8'hFD;
		16'h43AE: out_word = 8'h03;
		16'h43AF: out_word = 8'hCD;
		16'h43B0: out_word = 8'h80;
		16'h43B1: out_word = 8'h3D;
		16'h43B2: out_word = 8'hCD;
		16'h43B3: out_word = 8'h80;
		16'h43B4: out_word = 8'h3D;
		16'h43B5: out_word = 8'hED;
		16'h43B6: out_word = 8'h4B;
		16'h43B7: out_word = 8'h0A;
		16'h43B8: out_word = 8'h5E;
		16'h43B9: out_word = 8'hCD;
		16'h43BA: out_word = 8'hA9;
		16'h43BB: out_word = 8'h1D;
		16'h43BC: out_word = 8'h21;
		16'h43BD: out_word = 8'hD2;
		16'h43BE: out_word = 8'h29;
		16'h43BF: out_word = 8'hDF;
		16'h43C0: out_word = 8'hC3;
		16'h43C1: out_word = 8'hD3;
		16'h43C2: out_word = 8'h01;
		16'h43C3: out_word = 8'hF5;
		16'h43C4: out_word = 8'h3A;
		16'h43C5: out_word = 8'h0E;
		16'h43C6: out_word = 8'h5D;
		16'h43C7: out_word = 8'hFE;
		16'h43C8: out_word = 8'hFE;
		16'h43C9: out_word = 8'h20;
		16'h43CA: out_word = 8'h02;
		16'h43CB: out_word = 8'hF1;
		16'h43CC: out_word = 8'hC9;
		16'h43CD: out_word = 8'hF1;
		16'h43CE: out_word = 8'h32;
		16'h43CF: out_word = 8'h0F;
		16'h43D0: out_word = 8'h5D;
		16'h43D1: out_word = 8'h3A;
		16'h43D2: out_word = 8'h15;
		16'h43D3: out_word = 8'h5D;
		16'h43D4: out_word = 8'hB7;
		16'h43D5: out_word = 8'hCC;
		16'h43D6: out_word = 8'h07;
		16'h43D7: out_word = 8'h27;
		16'h43D8: out_word = 8'hC9;
		16'h43D9: out_word = 8'h21;
		16'h43DA: out_word = 8'h28;
		16'h43DB: out_word = 8'h2A;
		16'h43DC: out_word = 8'h3E;
		16'h43DD: out_word = 8'h01;
		16'h43DE: out_word = 8'hC3;
		16'h43DF: out_word = 8'h4A;
		16'h43E0: out_word = 8'h1C;
		16'h43E1: out_word = 8'h21;
		16'h43E2: out_word = 8'h66;
		16'h43E3: out_word = 8'h27;
		16'h43E4: out_word = 8'hAF;
		16'h43E5: out_word = 8'hC3;
		16'h43E6: out_word = 8'h4A;
		16'h43E7: out_word = 8'h1C;
		16'h43E8: out_word = 8'hAF;
		16'h43E9: out_word = 8'h32;
		16'h43EA: out_word = 8'hCC;
		16'h43EB: out_word = 8'h5C;
		16'h43EC: out_word = 8'hED;
		16'h43ED: out_word = 8'h5B;
		16'h43EE: out_word = 8'hCC;
		16'h43EF: out_word = 8'h5C;
		16'h43F0: out_word = 8'h16;
		16'h43F1: out_word = 8'h00;
		16'h43F2: out_word = 8'hCD;
		16'h43F3: out_word = 8'h4A;
		16'h43F4: out_word = 8'h29;
		16'h43F5: out_word = 8'h21;
		16'h43F6: out_word = 8'h25;
		16'h43F7: out_word = 8'h5D;
		16'h43F8: out_word = 8'h06;
		16'h43F9: out_word = 8'h01;
		16'h43FA: out_word = 8'hC3;
		16'h43FB: out_word = 8'h3D;
		16'h43FC: out_word = 8'h1E;
		16'h43FD: out_word = 8'hCD;
		16'h43FE: out_word = 8'h4A;
		16'h43FF: out_word = 8'h29;
		16'h4400: out_word = 8'h11;
		16'h4401: out_word = 8'h08;
		16'h4402: out_word = 8'h00;
		16'h4403: out_word = 8'h18;
		16'h4404: out_word = 8'hED;
		16'h4405: out_word = 8'hCD;
		16'h4406: out_word = 8'hFD;
		16'h4407: out_word = 8'h03;
		16'h4408: out_word = 8'h3A;
		16'h4409: out_word = 8'h0C;
		16'h440A: out_word = 8'h5E;
		16'h440B: out_word = 8'hFE;
		16'h440C: out_word = 8'h10;
		16'h440D: out_word = 8'h28;
		16'h440E: out_word = 8'h06;
		16'h440F: out_word = 8'h21;
		16'h4410: out_word = 8'hE2;
		16'h4411: out_word = 8'h29;
		16'h4412: out_word = 8'hDF;
		16'h4413: out_word = 8'h18;
		16'h4414: out_word = 8'hAB;
		16'h4415: out_word = 8'hCD;
		16'h4416: out_word = 8'h11;
		16'h4417: out_word = 8'h3E;
		16'h4418: out_word = 8'hCB;
		16'h4419: out_word = 8'h86;
		16'h441A: out_word = 8'hCB;
		16'h441B: out_word = 8'h8E;
		16'h441C: out_word = 8'h3A;
		16'h441D: out_word = 8'h08;
		16'h441E: out_word = 8'h5E;
		16'h441F: out_word = 8'hCB;
		16'h4420: out_word = 8'h47;
		16'h4421: out_word = 8'h20;
		16'h4422: out_word = 8'h02;
		16'h4423: out_word = 8'hCB;
		16'h4424: out_word = 8'hC6;
		16'h4425: out_word = 8'hCB;
		16'h4426: out_word = 8'h5F;
		16'h4427: out_word = 8'hC0;
		16'h4428: out_word = 8'hCB;
		16'h4429: out_word = 8'hCE;
		16'h442A: out_word = 8'hC9;
		16'h442B: out_word = 8'h2A;
		16'h442C: out_word = 8'h11;
		16'h442D: out_word = 8'h5D;
		16'h442E: out_word = 8'h23;
		16'h442F: out_word = 8'h7E;
		16'h4430: out_word = 8'hFE;
		16'h4431: out_word = 8'h0D;
		16'h4432: out_word = 8'hC9;
		16'h4433: out_word = 8'hCD;
		16'h4434: out_word = 8'h2B;
		16'h4435: out_word = 8'h04;
		16'h4436: out_word = 8'h01;
		16'h4437: out_word = 8'h02;
		16'h4438: out_word = 8'h00;
		16'h4439: out_word = 8'hED;
		16'h443A: out_word = 8'h43;
		16'h443B: out_word = 8'hDB;
		16'h443C: out_word = 8'h5C;
		16'h443D: out_word = 8'h28;
		16'h443E: out_word = 8'h2B;
		16'h443F: out_word = 8'hFE;
		16'h4440: out_word = 8'h23;
		16'h4441: out_word = 8'h20;
		16'h4442: out_word = 8'h1A;
		16'h4443: out_word = 8'h22;
		16'h4444: out_word = 8'h5D;
		16'h4445: out_word = 8'h5C;
		16'h4446: out_word = 8'hCD;
		16'h4447: out_word = 8'h0B;
		16'h4448: out_word = 8'h1E;
		16'h4449: out_word = 8'hCD;
		16'h444A: out_word = 8'h8C;
		16'h444B: out_word = 8'h1D;
		16'h444C: out_word = 8'hFE;
		16'h444D: out_word = 8'h0D;
		16'h444E: out_word = 8'h28;
		16'h444F: out_word = 8'h1A;
		16'h4450: out_word = 8'hFE;
		16'h4451: out_word = 8'h2C;
		16'h4452: out_word = 8'hC2;
		16'h4453: out_word = 8'h1A;
		16'h4454: out_word = 8'h1D;
		16'h4455: out_word = 8'hCD;
		16'h4456: out_word = 8'h2A;
		16'h4457: out_word = 8'h1E;
		16'h4458: out_word = 8'hCD;
		16'h4459: out_word = 8'hBD;
		16'h445A: out_word = 8'h1D;
		16'h445B: out_word = 8'h18;
		16'h445C: out_word = 8'h03;
		16'h445D: out_word = 8'hCD;
		16'h445E: out_word = 8'hDF;
		16'h445F: out_word = 8'h1D;
		16'h4460: out_word = 8'hCD;
		16'h4461: out_word = 8'h75;
		16'h4462: out_word = 8'h1D;
		16'h4463: out_word = 8'hCD;
		16'h4464: out_word = 8'hB5;
		16'h4465: out_word = 8'h1D;
		16'h4466: out_word = 8'hEB;
		16'h4467: out_word = 8'hCD;
		16'h4468: out_word = 8'h81;
		16'h4469: out_word = 8'h1C;
		16'h446A: out_word = 8'hCD;
		16'h446B: out_word = 8'h75;
		16'h446C: out_word = 8'h1D;
		16'h446D: out_word = 8'h3A;
		16'h446E: out_word = 8'hF6;
		16'h446F: out_word = 8'h5C;
		16'h4470: out_word = 8'h32;
		16'h4471: out_word = 8'hF9;
		16'h4472: out_word = 8'h5C;
		16'h4473: out_word = 8'hCD;
		16'h4474: out_word = 8'h05;
		16'h4475: out_word = 8'h04;
		16'h4476: out_word = 8'h3A;
		16'h4477: out_word = 8'hDB;
		16'h4478: out_word = 8'h5C;
		16'h4479: out_word = 8'hFE;
		16'h447A: out_word = 8'h02;
		16'h447B: out_word = 8'hF5;
		16'h447C: out_word = 8'hCC;
		16'h447D: out_word = 8'h97;
		16'h447E: out_word = 8'h1D;
		16'h447F: out_word = 8'hF1;
		16'h4480: out_word = 8'hFE;
		16'h4481: out_word = 8'h11;
		16'h4482: out_word = 8'hD2;
		16'h4483: out_word = 8'h1A;
		16'h4484: out_word = 8'h1D;
		16'h4485: out_word = 8'hCD;
		16'h4486: out_word = 8'h84;
		16'h4487: out_word = 8'h1D;
		16'h4488: out_word = 8'h3E;
		16'h4489: out_word = 8'hFF;
		16'h448A: out_word = 8'h32;
		16'h448B: out_word = 8'hF8;
		16'h448C: out_word = 8'h5C;
		16'h448D: out_word = 8'h21;
		16'h448E: out_word = 8'hF7;
		16'h448F: out_word = 8'h29;
		16'h4490: out_word = 8'hDF;
		16'h4491: out_word = 8'h21;
		16'h4492: out_word = 8'h1A;
		16'h4493: out_word = 8'h5E;
		16'h4494: out_word = 8'hDF;
		16'h4495: out_word = 8'hCD;
		16'h4496: out_word = 8'h80;
		16'h4497: out_word = 8'h3D;
		16'h4498: out_word = 8'h3A;
		16'h4499: out_word = 8'h09;
		16'h449A: out_word = 8'h5E;
		16'h449B: out_word = 8'h21;
		16'h449C: out_word = 8'h19;
		16'h449D: out_word = 8'h5E;
		16'h449E: out_word = 8'h96;
		16'h449F: out_word = 8'hE5;
		16'h44A0: out_word = 8'hCD;
		16'h44A1: out_word = 8'hA3;
		16'h44A2: out_word = 8'h1D;
		16'h44A3: out_word = 8'h21;
		16'h44A4: out_word = 8'h2B;
		16'h44A5: out_word = 8'h2A;
		16'h44A6: out_word = 8'hDF;
		16'h44A7: out_word = 8'hE1;
		16'h44A8: out_word = 8'h4E;
		16'h44A9: out_word = 8'hCD;
		16'h44AA: out_word = 8'hA4;
		16'h44AB: out_word = 8'h1D;
		16'h44AC: out_word = 8'h21;
		16'h44AD: out_word = 8'h1D;
		16'h44AE: out_word = 8'h2A;
		16'h44AF: out_word = 8'hDF;
		16'h44B0: out_word = 8'hCD;
		16'h44B1: out_word = 8'hE8;
		16'h44B2: out_word = 8'h03;
		16'h44B3: out_word = 8'h21;
		16'h44B4: out_word = 8'h25;
		16'h44B5: out_word = 8'h5D;
		16'h44B6: out_word = 8'hCD;
		16'h44B7: out_word = 8'hF6;
		16'h44B8: out_word = 8'h04;
		16'h44B9: out_word = 8'hCD;
		16'h44BA: out_word = 8'h80;
		16'h44BB: out_word = 8'h3D;
		16'h44BC: out_word = 8'h3A;
		16'h44BD: out_word = 8'hF6;
		16'h44BE: out_word = 8'h5C;
		16'h44BF: out_word = 8'hC6;
		16'h44C0: out_word = 8'h41;
		16'h44C1: out_word = 8'hD7;
		16'h44C2: out_word = 8'h06;
		16'h44C3: out_word = 8'h02;
		16'h44C4: out_word = 8'hCD;
		16'h44C5: out_word = 8'hF6;
		16'h44C6: out_word = 8'h04;
		16'h44C7: out_word = 8'hC5;
		16'h44C8: out_word = 8'h3E;
		16'h44C9: out_word = 8'h3A;
		16'h44CA: out_word = 8'hD7;
		16'h44CB: out_word = 8'hE5;
		16'h44CC: out_word = 8'hCD;
		16'h44CD: out_word = 8'h38;
		16'h44CE: out_word = 8'h29;
		16'h44CF: out_word = 8'h01;
		16'h44D0: out_word = 8'h0D;
		16'h44D1: out_word = 8'h00;
		16'h44D2: out_word = 8'hE1;
		16'h44D3: out_word = 8'hE5;
		16'h44D4: out_word = 8'h09;
		16'h44D5: out_word = 8'h4E;
		16'h44D6: out_word = 8'hC5;
		16'h44D7: out_word = 8'h79;
		16'h44D8: out_word = 8'h06;
		16'h44D9: out_word = 8'h02;
		16'h44DA: out_word = 8'hFE;
		16'h44DB: out_word = 8'h0A;
		16'h44DC: out_word = 8'h38;
		16'h44DD: out_word = 8'h01;
		16'h44DE: out_word = 8'h05;
		16'h44DF: out_word = 8'hFE;
		16'h44E0: out_word = 8'h64;
		16'h44E1: out_word = 8'h30;
		16'h44E2: out_word = 8'h05;
		16'h44E3: out_word = 8'h3E;
		16'h44E4: out_word = 8'h20;
		16'h44E5: out_word = 8'hD7;
		16'h44E6: out_word = 8'h10;
		16'h44E7: out_word = 8'hFB;
		16'h44E8: out_word = 8'hC1;
		16'h44E9: out_word = 8'hCD;
		16'h44EA: out_word = 8'hA9;
		16'h44EB: out_word = 8'h1D;
		16'h44EC: out_word = 8'hE1;
		16'h44ED: out_word = 8'hC1;
		16'h44EE: out_word = 8'h11;
		16'h44EF: out_word = 8'h10;
		16'h44F0: out_word = 8'h00;
		16'h44F1: out_word = 8'h19;
		16'h44F2: out_word = 8'h10;
		16'h44F3: out_word = 8'hD0;
		16'h44F4: out_word = 8'h18;
		16'h44F5: out_word = 8'hC0;
		16'h44F6: out_word = 8'hE5;
		16'h44F7: out_word = 8'hC5;
		16'h44F8: out_word = 8'h3A;
		16'h44F9: out_word = 8'hF9;
		16'h44FA: out_word = 8'h5C;
		16'h44FB: out_word = 8'h21;
		16'h44FC: out_word = 8'hF6;
		16'h44FD: out_word = 8'h5C;
		16'h44FE: out_word = 8'hBE;
		16'h44FF: out_word = 8'hC4;
		16'h4500: out_word = 8'hCB;
		16'h4501: out_word = 8'h3D;
		16'h4502: out_word = 8'hC1;
		16'h4503: out_word = 8'hE1;
		16'h4504: out_word = 8'hC3;
		16'h4505: out_word = 8'hC6;
		16'h4506: out_word = 8'h2F;
		16'h4507: out_word = 8'h11;
		16'h4508: out_word = 8'h10;
		16'h4509: out_word = 8'h00;
		16'h450A: out_word = 8'h19;
		16'h450B: out_word = 8'hC9;
		16'h450C: out_word = 8'hE5;
		16'h450D: out_word = 8'hC5;
		16'h450E: out_word = 8'h01;
		16'h450F: out_word = 8'hDB;
		16'h4510: out_word = 8'hA1;
		16'h4511: out_word = 8'h09;
		16'h4512: out_word = 8'h38;
		16'h4513: out_word = 8'h03;
		16'h4514: out_word = 8'hC1;
		16'h4515: out_word = 8'hE1;
		16'h4516: out_word = 8'hC9;
		16'h4517: out_word = 8'h21;
		16'h4518: out_word = 8'hCC;
		16'h4519: out_word = 8'h5C;
		16'h451A: out_word = 8'h34;
		16'h451B: out_word = 8'hCD;
		16'h451C: out_word = 8'hEC;
		16'h451D: out_word = 8'h03;
		16'h451E: out_word = 8'hC1;
		16'h451F: out_word = 8'hE1;
		16'h4520: out_word = 8'h21;
		16'h4521: out_word = 8'h25;
		16'h4522: out_word = 8'h5D;
		16'h4523: out_word = 8'hC9;
		16'h4524: out_word = 8'hE6;
		16'h4525: out_word = 8'hDF;
		16'h4526: out_word = 8'hDE;
		16'h4527: out_word = 8'h41;
		16'h4528: out_word = 8'hDA;
		16'h4529: out_word = 8'h1A;
		16'h452A: out_word = 8'h1D;
		16'h452B: out_word = 8'hFE;
		16'h452C: out_word = 8'h04;
		16'h452D: out_word = 8'hD2;
		16'h452E: out_word = 8'h1A;
		16'h452F: out_word = 8'h1D;
		16'h4530: out_word = 8'hC9;
		16'h4531: out_word = 8'hCD;
		16'h4532: out_word = 8'hB5;
		16'h4533: out_word = 8'h1D;
		16'h4534: out_word = 8'h79;
		16'h4535: out_word = 8'hB8;
		16'h4536: out_word = 8'hCA;
		16'h4537: out_word = 8'h1A;
		16'h4538: out_word = 8'h1D;
		16'h4539: out_word = 8'hC9;
		16'h453A: out_word = 8'hC3;
		16'h453B: out_word = 8'hD8;
		16'h453C: out_word = 8'h37;
		16'h453D: out_word = 8'hCD;
		16'h453E: out_word = 8'h75;
		16'h453F: out_word = 8'h1D;
		16'h4540: out_word = 8'hCD;
		16'h4541: out_word = 8'h2E;
		16'h4542: out_word = 8'h10;
		16'h4543: out_word = 8'hCD;
		16'h4544: out_word = 8'hB0;
		16'h4545: out_word = 8'h1C;
		16'h4546: out_word = 8'h3A;
		16'h4547: out_word = 8'hF6;
		16'h4548: out_word = 8'h5C;
		16'h4549: out_word = 8'h32;
		16'h454A: out_word = 8'hF8;
		16'h454B: out_word = 8'h5C;
		16'h454C: out_word = 8'hC2;
		16'h454D: out_word = 8'hD9;
		16'h454E: out_word = 8'h03;
		16'h454F: out_word = 8'hC5;
		16'h4550: out_word = 8'hCD;
		16'h4551: out_word = 8'h5D;
		16'h4552: out_word = 8'h16;
		16'h4553: out_word = 8'hCD;
		16'h4554: out_word = 8'hB0;
		16'h4555: out_word = 8'h1C;
		16'h4556: out_word = 8'hF5;
		16'h4557: out_word = 8'h3A;
		16'h4558: out_word = 8'hF8;
		16'h4559: out_word = 8'h5C;
		16'h455A: out_word = 8'h21;
		16'h455B: out_word = 8'hF6;
		16'h455C: out_word = 8'h5C;
		16'h455D: out_word = 8'hBE;
		16'h455E: out_word = 8'hC2;
		16'h455F: out_word = 8'h1A;
		16'h4560: out_word = 8'h1D;
		16'h4561: out_word = 8'hCD;
		16'h4562: out_word = 8'h05;
		16'h4563: out_word = 8'h04;
		16'h4564: out_word = 8'hF1;
		16'h4565: out_word = 8'hCA;
		16'h4566: out_word = 8'h50;
		16'h4567: out_word = 8'h1C;
		16'h4568: out_word = 8'hC1;
		16'h4569: out_word = 8'hCD;
		16'h456A: out_word = 8'h6B;
		16'h456B: out_word = 8'h16;
		16'h456C: out_word = 8'hCD;
		16'h456D: out_word = 8'h43;
		16'h456E: out_word = 8'h1E;
		16'h456F: out_word = 8'hC3;
		16'h4570: out_word = 8'hE1;
		16'h4571: out_word = 8'h03;
		16'h4572: out_word = 8'h3A;
		16'h4573: out_word = 8'h10;
		16'h4574: out_word = 8'h5D;
		16'h4575: out_word = 8'hB7;
		16'h4576: out_word = 8'hC9;
		16'h4577: out_word = 8'h3A;
		16'h4578: out_word = 8'h07;
		16'h4579: out_word = 8'h5D;
		16'h457A: out_word = 8'hB7;
		16'h457B: out_word = 8'hCA;
		16'h457C: out_word = 8'hD9;
		16'h457D: out_word = 8'h03;
		16'h457E: out_word = 8'hC3;
		16'h457F: out_word = 8'hE1;
		16'h4580: out_word = 8'h03;
		16'h4581: out_word = 8'hC5;
		16'h4582: out_word = 8'hCD;
		16'h4583: out_word = 8'h97;
		16'h4584: out_word = 8'h1D;
		16'h4585: out_word = 8'h3A;
		16'h4586: out_word = 8'hF6;
		16'h4587: out_word = 8'h5C;
		16'h4588: out_word = 8'hC6;
		16'h4589: out_word = 8'h41;
		16'h458A: out_word = 8'hCD;
		16'h458B: out_word = 8'h82;
		16'h458C: out_word = 8'h3D;
		16'h458D: out_word = 8'h3E;
		16'h458E: out_word = 8'h3A;
		16'h458F: out_word = 8'hCD;
		16'h4590: out_word = 8'h82;
		16'h4591: out_word = 8'h3D;
		16'h4592: out_word = 8'h21;
		16'h4593: out_word = 8'hDD;
		16'h4594: out_word = 8'h5C;
		16'h4595: out_word = 8'hCD;
		16'h4596: out_word = 8'h38;
		16'h4597: out_word = 8'h29;
		16'h4598: out_word = 8'h21;
		16'h4599: out_word = 8'h20;
		16'h459A: out_word = 8'h28;
		16'h459B: out_word = 8'hCD;
		16'h459C: out_word = 8'h07;
		16'h459D: out_word = 8'h27;
		16'h459E: out_word = 8'hCD;
		16'h459F: out_word = 8'h52;
		16'h45A0: out_word = 8'h10;
		16'h45A1: out_word = 8'hFE;
		16'h45A2: out_word = 8'h59;
		16'h45A3: out_word = 8'hF5;
		16'h45A4: out_word = 8'hCD;
		16'h45A5: out_word = 8'h97;
		16'h45A6: out_word = 8'h1D;
		16'h45A7: out_word = 8'hF1;
		16'h45A8: out_word = 8'hC1;
		16'h45A9: out_word = 8'hC0;
		16'h45AA: out_word = 8'hC5;
		16'h45AB: out_word = 8'hCD;
		16'h45AC: out_word = 8'h97;
		16'h45AD: out_word = 8'h1D;
		16'h45AE: out_word = 8'hC1;
		16'h45AF: out_word = 8'hCD;
		16'h45B0: out_word = 8'h81;
		16'h45B1: out_word = 8'h07;
		16'h45B2: out_word = 8'hAF;
		16'h45B3: out_word = 8'hC9;
		16'h45B4: out_word = 8'h3A;
		16'h45B5: out_word = 8'hE5;
		16'h45B6: out_word = 8'h5C;
		16'h45B7: out_word = 8'hFE;
		16'h45B8: out_word = 8'h23;
		16'h45B9: out_word = 8'h28;
		16'h45BA: out_word = 8'h02;
		16'h45BB: out_word = 8'hAF;
		16'h45BC: out_word = 8'hC9;
		16'h45BD: out_word = 8'h3E;
		16'h45BE: out_word = 8'h0A;
		16'h45BF: out_word = 8'h32;
		16'h45C0: out_word = 8'h06;
		16'h45C1: out_word = 8'h5D;
		16'h45C2: out_word = 8'hCD;
		16'h45C3: out_word = 8'hB3;
		16'h45C4: out_word = 8'h1C;
		16'h45C5: out_word = 8'h3E;
		16'h45C6: out_word = 8'h09;
		16'h45C7: out_word = 8'h32;
		16'h45C8: out_word = 8'h06;
		16'h45C9: out_word = 8'h5D;
		16'h45CA: out_word = 8'hC9;
		16'h45CB: out_word = 8'h3A;
		16'h45CC: out_word = 8'hDD;
		16'h45CD: out_word = 8'h5C;
		16'h45CE: out_word = 8'hFE;
		16'h45CF: out_word = 8'h2A;
		16'h45D0: out_word = 8'hC2;
		16'h45D1: out_word = 8'hD9;
		16'h45D2: out_word = 8'h03;
		16'h45D3: out_word = 8'hCD;
		16'h45D4: out_word = 8'hB5;
		16'h45D5: out_word = 8'h1D;
		16'h45D6: out_word = 8'hEB;
		16'h45D7: out_word = 8'hCD;
		16'h45D8: out_word = 8'h81;
		16'h45D9: out_word = 8'h1C;
		16'h45DA: out_word = 8'h7E;
		16'h45DB: out_word = 8'hFE;
		16'h45DC: out_word = 8'h2A;
		16'h45DD: out_word = 8'hC2;
		16'h45DE: out_word = 8'h1A;
		16'h45DF: out_word = 8'h1D;
		16'h45E0: out_word = 8'h3A;
		16'h45E1: out_word = 8'hF6;
		16'h45E2: out_word = 8'h5C;
		16'h45E3: out_word = 8'h32;
		16'h45E4: out_word = 8'hF9;
		16'h45E5: out_word = 8'h5C;
		16'h45E6: out_word = 8'h3A;
		16'h45E7: out_word = 8'hF9;
		16'h45E8: out_word = 8'h5C;
		16'h45E9: out_word = 8'hCD;
		16'h45EA: out_word = 8'hCB;
		16'h45EB: out_word = 8'h3D;
		16'h45EC: out_word = 8'hCD;
		16'h45ED: out_word = 8'h05;
		16'h45EE: out_word = 8'h04;
		16'h45EF: out_word = 8'h3E;
		16'h45F0: out_word = 8'hFF;
		16'h45F1: out_word = 8'h32;
		16'h45F2: out_word = 8'h0D;
		16'h45F3: out_word = 8'h5D;
		16'h45F4: out_word = 8'h3A;
		16'h45F5: out_word = 8'hF8;
		16'h45F6: out_word = 8'h5C;
		16'h45F7: out_word = 8'hCD;
		16'h45F8: out_word = 8'hCB;
		16'h45F9: out_word = 8'h3D;
		16'h45FA: out_word = 8'hCD;
		16'h45FB: out_word = 8'h05;
		16'h45FC: out_word = 8'h04;
		16'h45FD: out_word = 8'h3A;
		16'h45FE: out_word = 8'h0D;
		16'h45FF: out_word = 8'h5D;
		16'h4600: out_word = 8'h3C;
		16'h4601: out_word = 8'h32;
		16'h4602: out_word = 8'h0D;
		16'h4603: out_word = 8'h5D;
		16'h4604: out_word = 8'h4F;
		16'h4605: out_word = 8'hCD;
		16'h4606: out_word = 8'h5D;
		16'h4607: out_word = 8'h16;
		16'h4608: out_word = 8'h3A;
		16'h4609: out_word = 8'hDD;
		16'h460A: out_word = 8'h5C;
		16'h460B: out_word = 8'hFE;
		16'h460C: out_word = 8'h00;
		16'h460D: out_word = 8'hCA;
		16'h460E: out_word = 8'hE1;
		16'h460F: out_word = 8'h03;
		16'h4610: out_word = 8'hFE;
		16'h4611: out_word = 8'h01;
		16'h4612: out_word = 8'h28;
		16'h4613: out_word = 8'hE0;
		16'h4614: out_word = 8'h21;
		16'h4615: out_word = 8'hE6;
		16'h4616: out_word = 8'h5C;
		16'h4617: out_word = 8'h11;
		16'h4618: out_word = 8'hED;
		16'h4619: out_word = 8'h5C;
		16'h461A: out_word = 8'h01;
		16'h461B: out_word = 8'h07;
		16'h461C: out_word = 8'h00;
		16'h461D: out_word = 8'hED;
		16'h461E: out_word = 8'hB0;
		16'h461F: out_word = 8'h3A;
		16'h4620: out_word = 8'hF9;
		16'h4621: out_word = 8'h5C;
		16'h4622: out_word = 8'hCD;
		16'h4623: out_word = 8'hCB;
		16'h4624: out_word = 8'h3D;
		16'h4625: out_word = 8'hCD;
		16'h4626: out_word = 8'hB3;
		16'h4627: out_word = 8'h1C;
		16'h4628: out_word = 8'h20;
		16'h4629: out_word = 8'h0A;
		16'h462A: out_word = 8'hCD;
		16'h462B: out_word = 8'hB4;
		16'h462C: out_word = 8'h05;
		16'h462D: out_word = 8'h20;
		16'h462E: out_word = 8'h05;
		16'h462F: out_word = 8'hCD;
		16'h4630: out_word = 8'h81;
		16'h4631: out_word = 8'h05;
		16'h4632: out_word = 8'h20;
		16'h4633: out_word = 8'hC0;
		16'h4634: out_word = 8'hCD;
		16'h4635: out_word = 8'h3C;
		16'h4636: out_word = 8'h06;
		16'h4637: out_word = 8'hCD;
		16'h4638: out_word = 8'h43;
		16'h4639: out_word = 8'h1E;
		16'h463A: out_word = 8'h18;
		16'h463B: out_word = 8'hB8;
		16'h463C: out_word = 8'hCD;
		16'h463D: out_word = 8'hFD;
		16'h463E: out_word = 8'h03;
		16'h463F: out_word = 8'h3A;
		16'h4640: out_word = 8'h09;
		16'h4641: out_word = 8'h5E;
		16'h4642: out_word = 8'hFE;
		16'h4643: out_word = 8'h80;
		16'h4644: out_word = 8'hCA;
		16'h4645: out_word = 8'h23;
		16'h4646: out_word = 8'h27;
		16'h4647: out_word = 8'h21;
		16'h4648: out_word = 8'hED;
		16'h4649: out_word = 8'h5C;
		16'h464A: out_word = 8'h11;
		16'h464B: out_word = 8'hE6;
		16'h464C: out_word = 8'h5C;
		16'h464D: out_word = 8'h01;
		16'h464E: out_word = 8'h07;
		16'h464F: out_word = 8'h00;
		16'h4650: out_word = 8'hED;
		16'h4651: out_word = 8'hB0;
		16'h4652: out_word = 8'hED;
		16'h4653: out_word = 8'h5B;
		16'h4654: out_word = 8'hEA;
		16'h4655: out_word = 8'h5C;
		16'h4656: out_word = 8'h16;
		16'h4657: out_word = 8'h00;
		16'h4658: out_word = 8'hB7;
		16'h4659: out_word = 8'h2A;
		16'h465A: out_word = 8'h0A;
		16'h465B: out_word = 8'h5E;
		16'h465C: out_word = 8'hED;
		16'h465D: out_word = 8'h52;
		16'h465E: out_word = 8'hDA;
		16'h465F: out_word = 8'h45;
		16'h4660: out_word = 8'h1C;
		16'h4661: out_word = 8'h22;
		16'h4662: out_word = 8'h0A;
		16'h4663: out_word = 8'h5E;
		16'h4664: out_word = 8'h2A;
		16'h4665: out_word = 8'h06;
		16'h4666: out_word = 8'h5E;
		16'h4667: out_word = 8'h22;
		16'h4668: out_word = 8'hEB;
		16'h4669: out_word = 8'h5C;
		16'h466A: out_word = 8'hE5;
		16'h466B: out_word = 8'hCD;
		16'h466C: out_word = 8'h2F;
		16'h466D: out_word = 8'h07;
		16'h466E: out_word = 8'hE1;
		16'h466F: out_word = 8'h22;
		16'h4670: out_word = 8'hEB;
		16'h4671: out_word = 8'h5C;
		16'h4672: out_word = 8'h2A;
		16'h4673: out_word = 8'hF4;
		16'h4674: out_word = 8'h5C;
		16'h4675: out_word = 8'h22;
		16'h4676: out_word = 8'h06;
		16'h4677: out_word = 8'h5E;
		16'h4678: out_word = 8'h21;
		16'h4679: out_word = 8'h09;
		16'h467A: out_word = 8'h5E;
		16'h467B: out_word = 8'h34;
		16'h467C: out_word = 8'h4E;
		16'h467D: out_word = 8'h0D;
		16'h467E: out_word = 8'h06;
		16'h467F: out_word = 8'h00;
		16'h4680: out_word = 8'hC5;
		16'h4681: out_word = 8'h11;
		16'h4682: out_word = 8'h09;
		16'h4683: out_word = 8'h00;
		16'h4684: out_word = 8'hED;
		16'h4685: out_word = 8'h53;
		16'h4686: out_word = 8'hF4;
		16'h4687: out_word = 8'h5C;
		16'h4688: out_word = 8'hCD;
		16'h4689: out_word = 8'h43;
		16'h468A: out_word = 8'h1E;
		16'h468B: out_word = 8'hC1;
		16'h468C: out_word = 8'hCD;
		16'h468D: out_word = 8'h6B;
		16'h468E: out_word = 8'h16;
		16'h468F: out_word = 8'hC9;
		16'h4690: out_word = 8'h2A;
		16'h4691: out_word = 8'h11;
		16'h4692: out_word = 8'h5D;
		16'h4693: out_word = 8'h23;
		16'h4694: out_word = 8'h7E;
		16'h4695: out_word = 8'hE6;
		16'h4696: out_word = 8'hDF;
		16'h4697: out_word = 8'hFE;
		16'h4698: out_word = 8'h53;
		16'h4699: out_word = 8'hCA;
		16'h469A: out_word = 8'h60;
		16'h469B: out_word = 8'h13;
		16'h469C: out_word = 8'hFE;
		16'h469D: out_word = 8'h42;
		16'h469E: out_word = 8'hCA;
		16'h469F: out_word = 8'h2C;
		16'h46A0: out_word = 8'h15;
		16'h46A1: out_word = 8'hCD;
		16'h46A2: out_word = 8'hCD;
		16'h46A3: out_word = 8'h1D;
		16'h46A4: out_word = 8'hCD;
		16'h46A5: out_word = 8'h75;
		16'h46A6: out_word = 8'h1D;
		16'h46A7: out_word = 8'hCD;
		16'h46A8: out_word = 8'h6F;
		16'h46A9: out_word = 8'h16;
		16'h46AA: out_word = 8'hCD;
		16'h46AB: out_word = 8'h2E;
		16'h46AC: out_word = 8'h10;
		16'h46AD: out_word = 8'hCD;
		16'h46AE: out_word = 8'hB0;
		16'h46AF: out_word = 8'h1C;
		16'h46B0: out_word = 8'h3A;
		16'h46B1: out_word = 8'hF6;
		16'h46B2: out_word = 8'h5C;
		16'h46B3: out_word = 8'h32;
		16'h46B4: out_word = 8'hF8;
		16'h46B5: out_word = 8'h5C;
		16'h46B6: out_word = 8'hC2;
		16'h46B7: out_word = 8'hCB;
		16'h46B8: out_word = 8'h05;
		16'h46B9: out_word = 8'hCD;
		16'h46BA: out_word = 8'h5D;
		16'h46BB: out_word = 8'h16;
		16'h46BC: out_word = 8'h21;
		16'h46BD: out_word = 8'hE6;
		16'h46BE: out_word = 8'h5C;
		16'h46BF: out_word = 8'h11;
		16'h46C0: out_word = 8'hED;
		16'h46C1: out_word = 8'h5C;
		16'h46C2: out_word = 8'h01;
		16'h46C3: out_word = 8'h07;
		16'h46C4: out_word = 8'h00;
		16'h46C5: out_word = 8'hED;
		16'h46C6: out_word = 8'hB0;
		16'h46C7: out_word = 8'hCD;
		16'h46C8: out_word = 8'hB0;
		16'h46C9: out_word = 8'h1C;
		16'h46CA: out_word = 8'hF5;
		16'h46CB: out_word = 8'hC5;
		16'h46CC: out_word = 8'h3A;
		16'h46CD: out_word = 8'hF6;
		16'h46CE: out_word = 8'h5C;
		16'h46CF: out_word = 8'h32;
		16'h46D0: out_word = 8'hF9;
		16'h46D1: out_word = 8'h5C;
		16'h46D2: out_word = 8'h3A;
		16'h46D3: out_word = 8'hF8;
		16'h46D4: out_word = 8'h5C;
		16'h46D5: out_word = 8'hCD;
		16'h46D6: out_word = 8'hCB;
		16'h46D7: out_word = 8'h3D;
		16'h46D8: out_word = 8'hCD;
		16'h46D9: out_word = 8'h05;
		16'h46DA: out_word = 8'h04;
		16'h46DB: out_word = 8'h3A;
		16'h46DC: out_word = 8'hF9;
		16'h46DD: out_word = 8'h5C;
		16'h46DE: out_word = 8'hCD;
		16'h46DF: out_word = 8'hCB;
		16'h46E0: out_word = 8'h3D;
		16'h46E1: out_word = 8'hCD;
		16'h46E2: out_word = 8'h05;
		16'h46E3: out_word = 8'h04;
		16'h46E4: out_word = 8'hC1;
		16'h46E5: out_word = 8'hF1;
		16'h46E6: out_word = 8'h20;
		16'h46E7: out_word = 8'h0B;
		16'h46E8: out_word = 8'hCD;
		16'h46E9: out_word = 8'hB4;
		16'h46EA: out_word = 8'h05;
		16'h46EB: out_word = 8'h20;
		16'h46EC: out_word = 8'h06;
		16'h46ED: out_word = 8'hCD;
		16'h46EE: out_word = 8'h81;
		16'h46EF: out_word = 8'h05;
		16'h46F0: out_word = 8'hC2;
		16'h46F1: out_word = 8'hE1;
		16'h46F2: out_word = 8'h03;
		16'h46F3: out_word = 8'hCD;
		16'h46F4: out_word = 8'h3C;
		16'h46F5: out_word = 8'h06;
		16'h46F6: out_word = 8'hCD;
		16'h46F7: out_word = 8'h43;
		16'h46F8: out_word = 8'h1E;
		16'h46F9: out_word = 8'h3A;
		16'h46FA: out_word = 8'hE5;
		16'h46FB: out_word = 8'h5C;
		16'h46FC: out_word = 8'hFE;
		16'h46FD: out_word = 8'h23;
		16'h46FE: out_word = 8'hC2;
		16'h46FF: out_word = 8'hE1;
		16'h4700: out_word = 8'h03;
		16'h4701: out_word = 8'h3E;
		16'h4702: out_word = 8'h0A;
		16'h4703: out_word = 8'h32;
		16'h4704: out_word = 8'h06;
		16'h4705: out_word = 8'h5D;
		16'h4706: out_word = 8'h21;
		16'h4707: out_word = 8'hE6;
		16'h4708: out_word = 8'h5C;
		16'h4709: out_word = 8'h34;
		16'h470A: out_word = 8'h3A;
		16'h470B: out_word = 8'hF8;
		16'h470C: out_word = 8'h5C;
		16'h470D: out_word = 8'hCD;
		16'h470E: out_word = 8'hCB;
		16'h470F: out_word = 8'h3D;
		16'h4710: out_word = 8'hCD;
		16'h4711: out_word = 8'hB4;
		16'h4712: out_word = 8'h05;
		16'h4713: out_word = 8'hC2;
		16'h4714: out_word = 8'hE1;
		16'h4715: out_word = 8'h03;
		16'h4716: out_word = 8'hCD;
		16'h4717: out_word = 8'h5D;
		16'h4718: out_word = 8'h16;
		16'h4719: out_word = 8'h21;
		16'h471A: out_word = 8'hE6;
		16'h471B: out_word = 8'h5C;
		16'h471C: out_word = 8'h11;
		16'h471D: out_word = 8'hED;
		16'h471E: out_word = 8'h5C;
		16'h471F: out_word = 8'h01;
		16'h4720: out_word = 8'h07;
		16'h4721: out_word = 8'h00;
		16'h4722: out_word = 8'hED;
		16'h4723: out_word = 8'hB0;
		16'h4724: out_word = 8'h3A;
		16'h4725: out_word = 8'hF9;
		16'h4726: out_word = 8'h5C;
		16'h4727: out_word = 8'hCD;
		16'h4728: out_word = 8'hCB;
		16'h4729: out_word = 8'h3D;
		16'h472A: out_word = 8'hCD;
		16'h472B: out_word = 8'h05;
		16'h472C: out_word = 8'h04;
		16'h472D: out_word = 8'h18;
		16'h472E: out_word = 8'hC4;
		16'h472F: out_word = 8'h3A;
		16'h4730: out_word = 8'hF1;
		16'h4731: out_word = 8'h5C;
		16'h4732: out_word = 8'hB7;
		16'h4733: out_word = 8'hC8;
		16'h4734: out_word = 8'hE5;
		16'h4735: out_word = 8'h21;
		16'h4736: out_word = 8'h23;
		16'h4737: out_word = 8'h5D;
		16'h4738: out_word = 8'h96;
		16'h4739: out_word = 8'hE1;
		16'h473A: out_word = 8'h30;
		16'h473B: out_word = 8'h39;
		16'h473C: out_word = 8'h3A;
		16'h473D: out_word = 8'hF1;
		16'h473E: out_word = 8'h5C;
		16'h473F: out_word = 8'h47;
		16'h4740: out_word = 8'hAF;
		16'h4741: out_word = 8'h32;
		16'h4742: out_word = 8'hF1;
		16'h4743: out_word = 8'h5C;
		16'h4744: out_word = 8'hC5;
		16'h4745: out_word = 8'h3A;
		16'h4746: out_word = 8'hF8;
		16'h4747: out_word = 8'h5C;
		16'h4748: out_word = 8'hCD;
		16'h4749: out_word = 8'hCB;
		16'h474A: out_word = 8'h3D;
		16'h474B: out_word = 8'hC1;
		16'h474C: out_word = 8'hC5;
		16'h474D: out_word = 8'h2A;
		16'h474E: out_word = 8'hCF;
		16'h474F: out_word = 8'h5C;
		16'h4750: out_word = 8'hE5;
		16'h4751: out_word = 8'hED;
		16'h4752: out_word = 8'h5B;
		16'h4753: out_word = 8'hF2;
		16'h4754: out_word = 8'h5C;
		16'h4755: out_word = 8'hCD;
		16'h4756: out_word = 8'h3D;
		16'h4757: out_word = 8'h1E;
		16'h4758: out_word = 8'h2A;
		16'h4759: out_word = 8'hF4;
		16'h475A: out_word = 8'h5C;
		16'h475B: out_word = 8'h22;
		16'h475C: out_word = 8'hF2;
		16'h475D: out_word = 8'h5C;
		16'h475E: out_word = 8'h3A;
		16'h475F: out_word = 8'hF9;
		16'h4760: out_word = 8'h5C;
		16'h4761: out_word = 8'hCD;
		16'h4762: out_word = 8'hCB;
		16'h4763: out_word = 8'h3D;
		16'h4764: out_word = 8'hE1;
		16'h4765: out_word = 8'hC1;
		16'h4766: out_word = 8'hED;
		16'h4767: out_word = 8'h5B;
		16'h4768: out_word = 8'hEB;
		16'h4769: out_word = 8'h5C;
		16'h476A: out_word = 8'hCD;
		16'h476B: out_word = 8'h4D;
		16'h476C: out_word = 8'h1E;
		16'h476D: out_word = 8'h2A;
		16'h476E: out_word = 8'hF4;
		16'h476F: out_word = 8'h5C;
		16'h4770: out_word = 8'h22;
		16'h4771: out_word = 8'hEB;
		16'h4772: out_word = 8'h5C;
		16'h4773: out_word = 8'h18;
		16'h4774: out_word = 8'hBA;
		16'h4775: out_word = 8'h32;
		16'h4776: out_word = 8'hF1;
		16'h4777: out_word = 8'h5C;
		16'h4778: out_word = 8'hE5;
		16'h4779: out_word = 8'h21;
		16'h477A: out_word = 8'h23;
		16'h477B: out_word = 8'h5D;
		16'h477C: out_word = 8'h46;
		16'h477D: out_word = 8'hE1;
		16'h477E: out_word = 8'hAF;
		16'h477F: out_word = 8'h18;
		16'h4780: out_word = 8'hC3;
		16'h4781: out_word = 8'hAF;
		16'h4782: out_word = 8'h32;
		16'h4783: out_word = 8'h07;
		16'h4784: out_word = 8'h5D;
		16'h4785: out_word = 8'h18;
		16'h4786: out_word = 8'h19;
		16'h4787: out_word = 8'hCD;
		16'h4788: out_word = 8'hDF;
		16'h4789: out_word = 8'h1D;
		16'h478A: out_word = 8'hCD;
		16'h478B: out_word = 8'h75;
		16'h478C: out_word = 8'h1D;
		16'h478D: out_word = 8'hCD;
		16'h478E: out_word = 8'h2E;
		16'h478F: out_word = 8'h10;
		16'h4790: out_word = 8'hAF;
		16'h4791: out_word = 8'h32;
		16'h4792: out_word = 8'h07;
		16'h4793: out_word = 8'h5D;
		16'h4794: out_word = 8'hCD;
		16'h4795: out_word = 8'h2F;
		16'h4796: out_word = 8'h29;
		16'h4797: out_word = 8'hCD;
		16'h4798: out_word = 8'hA0;
		16'h4799: out_word = 8'h07;
		16'h479A: out_word = 8'hC2;
		16'h479B: out_word = 8'h77;
		16'h479C: out_word = 8'h05;
		16'h479D: out_word = 8'hC3;
		16'h479E: out_word = 8'hE1;
		16'h479F: out_word = 8'h03;
		16'h47A0: out_word = 8'h3A;
		16'h47A1: out_word = 8'hDD;
		16'h47A2: out_word = 8'h5C;
		16'h47A3: out_word = 8'h32;
		16'h47A4: out_word = 8'h08;
		16'h47A5: out_word = 8'h5D;
		16'h47A6: out_word = 8'hC0;
		16'h47A7: out_word = 8'h21;
		16'h47A8: out_word = 8'h07;
		16'h47A9: out_word = 8'h5D;
		16'h47AA: out_word = 8'h34;
		16'h47AB: out_word = 8'hC5;
		16'h47AC: out_word = 8'hCD;
		16'h47AD: out_word = 8'hFD;
		16'h47AE: out_word = 8'h03;
		16'h47AF: out_word = 8'h3A;
		16'h47B0: out_word = 8'h09;
		16'h47B1: out_word = 8'h5E;
		16'h47B2: out_word = 8'hC1;
		16'h47B3: out_word = 8'h0C;
		16'h47B4: out_word = 8'hB9;
		16'h47B5: out_word = 8'h20;
		16'h47B6: out_word = 8'h05;
		16'h47B7: out_word = 8'h3D;
		16'h47B8: out_word = 8'h32;
		16'h47B9: out_word = 8'h09;
		16'h47BA: out_word = 8'h5E;
		16'h47BB: out_word = 8'hAF;
		16'h47BC: out_word = 8'hF5;
		16'h47BD: out_word = 8'h28;
		16'h47BE: out_word = 8'h04;
		16'h47BF: out_word = 8'h21;
		16'h47C0: out_word = 8'h19;
		16'h47C1: out_word = 8'h5E;
		16'h47C2: out_word = 8'h34;
		16'h47C3: out_word = 8'hC5;
		16'h47C4: out_word = 8'hCD;
		16'h47C5: out_word = 8'h43;
		16'h47C6: out_word = 8'h1E;
		16'h47C7: out_word = 8'hC1;
		16'h47C8: out_word = 8'h0D;
		16'h47C9: out_word = 8'hCD;
		16'h47CA: out_word = 8'h5D;
		16'h47CB: out_word = 8'h16;
		16'h47CC: out_word = 8'hF1;
		16'h47CD: out_word = 8'hCA;
		16'h47CE: out_word = 8'hD2;
		16'h47CF: out_word = 8'h07;
		16'h47D0: out_word = 8'h3E;
		16'h47D1: out_word = 8'h01;
		16'h47D2: out_word = 8'h32;
		16'h47D3: out_word = 8'hDD;
		16'h47D4: out_word = 8'h5C;
		16'h47D5: out_word = 8'hF5;
		16'h47D6: out_word = 8'hCD;
		16'h47D7: out_word = 8'h40;
		16'h47D8: out_word = 8'h1E;
		16'h47D9: out_word = 8'h3A;
		16'h47DA: out_word = 8'h08;
		16'h47DB: out_word = 8'h5D;
		16'h47DC: out_word = 8'h32;
		16'h47DD: out_word = 8'hDD;
		16'h47DE: out_word = 8'h5C;
		16'h47DF: out_word = 8'hF1;
		16'h47E0: out_word = 8'h28;
		16'h47E1: out_word = 8'h05;
		16'h47E2: out_word = 8'hCD;
		16'h47E3: out_word = 8'hB3;
		16'h47E4: out_word = 8'h1C;
		16'h47E5: out_word = 8'h18;
		16'h47E6: out_word = 8'hB9;
		16'h47E7: out_word = 8'hCD;
		16'h47E8: out_word = 8'hFD;
		16'h47E9: out_word = 8'h03;
		16'h47EA: out_word = 8'h2A;
		16'h47EB: out_word = 8'hEB;
		16'h47EC: out_word = 8'h5C;
		16'h47ED: out_word = 8'h22;
		16'h47EE: out_word = 8'h06;
		16'h47EF: out_word = 8'h5E;
		16'h47F0: out_word = 8'hED;
		16'h47F1: out_word = 8'h5B;
		16'h47F2: out_word = 8'hEA;
		16'h47F3: out_word = 8'h5C;
		16'h47F4: out_word = 8'h2A;
		16'h47F5: out_word = 8'h0A;
		16'h47F6: out_word = 8'h5E;
		16'h47F7: out_word = 8'h16;
		16'h47F8: out_word = 8'h00;
		16'h47F9: out_word = 8'h19;
		16'h47FA: out_word = 8'h22;
		16'h47FB: out_word = 8'h0A;
		16'h47FC: out_word = 8'h5E;
		16'h47FD: out_word = 8'hC3;
		16'h47FE: out_word = 8'h43;
		16'h47FF: out_word = 8'h1E;
		16'h4800: out_word = 8'hE6;
		16'h4801: out_word = 8'hFC;
		16'h4802: out_word = 8'hC3;
		16'h4803: out_word = 8'h9A;
		16'h4804: out_word = 8'h3D;
		16'h4805: out_word = 8'hE5;
		16'h4806: out_word = 8'hC5;
		16'h4807: out_word = 8'hD5;
		16'h4808: out_word = 8'hF5;
		16'h4809: out_word = 8'hCD;
		16'h480A: out_word = 8'hF1;
		16'h480B: out_word = 8'h20;
		16'h480C: out_word = 8'hF1;
		16'h480D: out_word = 8'hCD;
		16'h480E: out_word = 8'h94;
		16'h480F: out_word = 8'h3D;
		16'h4810: out_word = 8'hCD;
		16'h4811: out_word = 8'hF1;
		16'h4812: out_word = 8'h20;
		16'h4813: out_word = 8'hD1;
		16'h4814: out_word = 8'hC1;
		16'h4815: out_word = 8'hE1;
		16'h4816: out_word = 8'hC9;
		16'h4817: out_word = 8'hE6;
		16'h4818: out_word = 8'h3F;
		16'h4819: out_word = 8'h6F;
		16'h481A: out_word = 8'h26;
		16'h481B: out_word = 8'h00;
		16'h481C: out_word = 8'h29;
		16'h481D: out_word = 8'h29;
		16'h481E: out_word = 8'h29;
		16'h481F: out_word = 8'h01;
		16'h4820: out_word = 8'h00;
		16'h4821: out_word = 8'h0C;
		16'h4822: out_word = 8'h09;
		16'h4823: out_word = 8'h11;
		16'h4824: out_word = 8'h92;
		16'h4825: out_word = 8'h5C;
		16'h4826: out_word = 8'h01;
		16'h4827: out_word = 8'h08;
		16'h4828: out_word = 8'h00;
		16'h4829: out_word = 8'hED;
		16'h482A: out_word = 8'hB0;
		16'h482B: out_word = 8'h3E;
		16'h482C: out_word = 8'hC9;
		16'h482D: out_word = 8'h32;
		16'h482E: out_word = 8'h9A;
		16'h482F: out_word = 8'h5C;
		16'h4830: out_word = 8'hC3;
		16'h4831: out_word = 8'h9A;
		16'h4832: out_word = 8'h5C;
		16'h4833: out_word = 8'h3A;
		16'h4834: out_word = 8'hF6;
		16'h4835: out_word = 8'h5C;
		16'h4836: out_word = 8'hFE;
		16'h4837: out_word = 8'h03;
		16'h4838: out_word = 8'h28;
		16'h4839: out_word = 8'h0E;
		16'h483A: out_word = 8'h3E;
		16'h483B: out_word = 8'h0D;
		16'h483C: out_word = 8'hD7;
		16'h483D: out_word = 8'h21;
		16'h483E: out_word = 8'h5E;
		16'h483F: out_word = 8'h33;
		16'h4840: out_word = 8'hDF;
		16'h4841: out_word = 8'hCD;
		16'h4842: out_word = 8'h52;
		16'h4843: out_word = 8'h10;
		16'h4844: out_word = 8'hFE;
		16'h4845: out_word = 8'h52;
		16'h4846: out_word = 8'h28;
		16'h4847: out_word = 8'h03;
		16'h4848: out_word = 8'hC3;
		16'h4849: out_word = 8'hD3;
		16'h484A: out_word = 8'h01;
		16'h484B: out_word = 8'hE7;
		16'h484C: out_word = 8'h6E;
		16'h484D: out_word = 8'h0D;
		16'h484E: out_word = 8'hE7;
		16'h484F: out_word = 8'h8E;
		16'h4850: out_word = 8'h02;
		16'h4851: out_word = 8'h20;
		16'h4852: out_word = 8'hFB;
		16'h4853: out_word = 8'hE7;
		16'h4854: out_word = 8'h1E;
		16'h4855: out_word = 8'h03;
		16'h4856: out_word = 8'h38;
		16'h4857: out_word = 8'hF6;
		16'h4858: out_word = 8'hC3;
		16'h4859: out_word = 8'hDD;
		16'h485A: out_word = 8'h1E;
		16'h485B: out_word = 8'hFF;
		16'h485C: out_word = 8'hFF;
		16'h485D: out_word = 8'hFF;
		16'h485E: out_word = 8'hFF;
		16'h485F: out_word = 8'hFF;
		16'h4860: out_word = 8'hFF;
		16'h4861: out_word = 8'hFF;
		16'h4862: out_word = 8'hFF;
		16'h4863: out_word = 8'hFF;
		16'h4864: out_word = 8'hFF;
		16'h4865: out_word = 8'hFF;
		16'h4866: out_word = 8'hFF;
		16'h4867: out_word = 8'hFF;
		16'h4868: out_word = 8'hFF;
		16'h4869: out_word = 8'hFF;
		16'h486A: out_word = 8'hFF;
		16'h486B: out_word = 8'hFF;
		16'h486C: out_word = 8'hFF;
		16'h486D: out_word = 8'hFF;
		16'h486E: out_word = 8'hFF;
		16'h486F: out_word = 8'hFF;
		16'h4870: out_word = 8'hFF;
		16'h4871: out_word = 8'hFF;
		16'h4872: out_word = 8'hFF;
		16'h4873: out_word = 8'hFF;
		16'h4874: out_word = 8'hFF;
		16'h4875: out_word = 8'hFF;
		16'h4876: out_word = 8'hFF;
		16'h4877: out_word = 8'hFF;
		16'h4878: out_word = 8'hFF;
		16'h4879: out_word = 8'hFF;
		16'h487A: out_word = 8'hFF;
		16'h487B: out_word = 8'hFF;
		16'h487C: out_word = 8'hFF;
		16'h487D: out_word = 8'hFF;
		16'h487E: out_word = 8'hFF;
		16'h487F: out_word = 8'hFF;
		16'h4880: out_word = 8'hFF;
		16'h4881: out_word = 8'hFF;
		16'h4882: out_word = 8'hFF;
		16'h4883: out_word = 8'hFF;
		16'h4884: out_word = 8'hFF;
		16'h4885: out_word = 8'hFF;
		16'h4886: out_word = 8'hFF;
		16'h4887: out_word = 8'hFF;
		16'h4888: out_word = 8'hFF;
		16'h4889: out_word = 8'hFF;
		16'h488A: out_word = 8'hFF;
		16'h488B: out_word = 8'hFF;
		16'h488C: out_word = 8'hFF;
		16'h488D: out_word = 8'hFF;
		16'h488E: out_word = 8'hFF;
		16'h488F: out_word = 8'hFF;
		16'h4890: out_word = 8'hFF;
		16'h4891: out_word = 8'hFF;
		16'h4892: out_word = 8'hFF;
		16'h4893: out_word = 8'hFF;
		16'h4894: out_word = 8'hFF;
		16'h4895: out_word = 8'hFF;
		16'h4896: out_word = 8'hFF;
		16'h4897: out_word = 8'hFF;
		16'h4898: out_word = 8'hFF;
		16'h4899: out_word = 8'hFF;
		16'h489A: out_word = 8'hFF;
		16'h489B: out_word = 8'hFF;
		16'h489C: out_word = 8'hFF;
		16'h489D: out_word = 8'hFF;
		16'h489E: out_word = 8'hFF;
		16'h489F: out_word = 8'hFF;
		16'h48A0: out_word = 8'hFF;
		16'h48A1: out_word = 8'hFF;
		16'h48A2: out_word = 8'hFF;
		16'h48A3: out_word = 8'hFF;
		16'h48A4: out_word = 8'hFF;
		16'h48A5: out_word = 8'hFF;
		16'h48A6: out_word = 8'hFF;
		16'h48A7: out_word = 8'hFF;
		16'h48A8: out_word = 8'hFF;
		16'h48A9: out_word = 8'hFF;
		16'h48AA: out_word = 8'hFF;
		16'h48AB: out_word = 8'hFF;
		16'h48AC: out_word = 8'hFF;
		16'h48AD: out_word = 8'hFF;
		16'h48AE: out_word = 8'hFF;
		16'h48AF: out_word = 8'hFF;
		16'h48B0: out_word = 8'hFF;
		16'h48B1: out_word = 8'hFF;
		16'h48B2: out_word = 8'hFF;
		16'h48B3: out_word = 8'hFF;
		16'h48B4: out_word = 8'hFF;
		16'h48B5: out_word = 8'hFF;
		16'h48B6: out_word = 8'hFF;
		16'h48B7: out_word = 8'hFF;
		16'h48B8: out_word = 8'hFF;
		16'h48B9: out_word = 8'hFF;
		16'h48BA: out_word = 8'hFF;
		16'h48BB: out_word = 8'hFF;
		16'h48BC: out_word = 8'hFF;
		16'h48BD: out_word = 8'hFF;
		16'h48BE: out_word = 8'hFF;
		16'h48BF: out_word = 8'hFF;
		16'h48C0: out_word = 8'hFF;
		16'h48C1: out_word = 8'hFF;
		16'h48C2: out_word = 8'hFF;
		16'h48C3: out_word = 8'hFF;
		16'h48C4: out_word = 8'hFF;
		16'h48C5: out_word = 8'hFF;
		16'h48C6: out_word = 8'hFF;
		16'h48C7: out_word = 8'hFF;
		16'h48C8: out_word = 8'hFF;
		16'h48C9: out_word = 8'hFF;
		16'h48CA: out_word = 8'hFF;
		16'h48CB: out_word = 8'hFF;
		16'h48CC: out_word = 8'hFF;
		16'h48CD: out_word = 8'hFF;
		16'h48CE: out_word = 8'hFF;
		16'h48CF: out_word = 8'hFF;
		16'h48D0: out_word = 8'hFF;
		16'h48D1: out_word = 8'hFF;
		16'h48D2: out_word = 8'hFF;
		16'h48D3: out_word = 8'hFF;
		16'h48D4: out_word = 8'hFF;
		16'h48D5: out_word = 8'hFF;
		16'h48D6: out_word = 8'hFF;
		16'h48D7: out_word = 8'hFF;
		16'h48D8: out_word = 8'hFF;
		16'h48D9: out_word = 8'hFF;
		16'h48DA: out_word = 8'hFF;
		16'h48DB: out_word = 8'hFF;
		16'h48DC: out_word = 8'hFF;
		16'h48DD: out_word = 8'hFF;
		16'h48DE: out_word = 8'hFF;
		16'h48DF: out_word = 8'hFF;
		16'h48E0: out_word = 8'hFF;
		16'h48E1: out_word = 8'hFF;
		16'h48E2: out_word = 8'hFF;
		16'h48E3: out_word = 8'hFF;
		16'h48E4: out_word = 8'hFF;
		16'h48E5: out_word = 8'hFF;
		16'h48E6: out_word = 8'hFF;
		16'h48E7: out_word = 8'hFF;
		16'h48E8: out_word = 8'hFF;
		16'h48E9: out_word = 8'hFF;
		16'h48EA: out_word = 8'hFF;
		16'h48EB: out_word = 8'hFF;
		16'h48EC: out_word = 8'hFF;
		16'h48ED: out_word = 8'hFF;
		16'h48EE: out_word = 8'hFF;
		16'h48EF: out_word = 8'hFF;
		16'h48F0: out_word = 8'hFF;
		16'h48F1: out_word = 8'hFF;
		16'h48F2: out_word = 8'hFF;
		16'h48F3: out_word = 8'hFF;
		16'h48F4: out_word = 8'hFF;
		16'h48F5: out_word = 8'hFF;
		16'h48F6: out_word = 8'hFF;
		16'h48F7: out_word = 8'hFF;
		16'h48F8: out_word = 8'hFF;
		16'h48F9: out_word = 8'hFF;
		16'h48FA: out_word = 8'hFF;
		16'h48FB: out_word = 8'hFF;
		16'h48FC: out_word = 8'hFF;
		16'h48FD: out_word = 8'hFF;
		16'h48FE: out_word = 8'hFF;
		16'h48FF: out_word = 8'hFF;
		16'h4900: out_word = 8'hFF;
		16'h4901: out_word = 8'hFF;
		16'h4902: out_word = 8'hFF;
		16'h4903: out_word = 8'hFF;
		16'h4904: out_word = 8'hFF;
		16'h4905: out_word = 8'hFF;
		16'h4906: out_word = 8'hFF;
		16'h4907: out_word = 8'hFF;
		16'h4908: out_word = 8'hFF;
		16'h4909: out_word = 8'hFF;
		16'h490A: out_word = 8'hFF;
		16'h490B: out_word = 8'hFF;
		16'h490C: out_word = 8'hFF;
		16'h490D: out_word = 8'hFF;
		16'h490E: out_word = 8'hFF;
		16'h490F: out_word = 8'hFF;
		16'h4910: out_word = 8'hFF;
		16'h4911: out_word = 8'hFF;
		16'h4912: out_word = 8'hFF;
		16'h4913: out_word = 8'hFF;
		16'h4914: out_word = 8'hFF;
		16'h4915: out_word = 8'hFF;
		16'h4916: out_word = 8'hFF;
		16'h4917: out_word = 8'hFF;
		16'h4918: out_word = 8'hFF;
		16'h4919: out_word = 8'hFF;
		16'h491A: out_word = 8'hFF;
		16'h491B: out_word = 8'hFF;
		16'h491C: out_word = 8'hFF;
		16'h491D: out_word = 8'hFF;
		16'h491E: out_word = 8'hFF;
		16'h491F: out_word = 8'hFF;
		16'h4920: out_word = 8'hFF;
		16'h4921: out_word = 8'hFF;
		16'h4922: out_word = 8'hFF;
		16'h4923: out_word = 8'hFF;
		16'h4924: out_word = 8'hFF;
		16'h4925: out_word = 8'hFF;
		16'h4926: out_word = 8'hFF;
		16'h4927: out_word = 8'hFF;
		16'h4928: out_word = 8'hFF;
		16'h4929: out_word = 8'hFF;
		16'h492A: out_word = 8'hFF;
		16'h492B: out_word = 8'hFF;
		16'h492C: out_word = 8'hFF;
		16'h492D: out_word = 8'hFF;
		16'h492E: out_word = 8'hFF;
		16'h492F: out_word = 8'hFF;
		16'h4930: out_word = 8'hFF;
		16'h4931: out_word = 8'hFF;
		16'h4932: out_word = 8'hFF;
		16'h4933: out_word = 8'hFF;
		16'h4934: out_word = 8'hFF;
		16'h4935: out_word = 8'hFF;
		16'h4936: out_word = 8'hFF;
		16'h4937: out_word = 8'hFF;
		16'h4938: out_word = 8'hFF;
		16'h4939: out_word = 8'hFF;
		16'h493A: out_word = 8'hFF;
		16'h493B: out_word = 8'hFF;
		16'h493C: out_word = 8'hFF;
		16'h493D: out_word = 8'hFF;
		16'h493E: out_word = 8'hFF;
		16'h493F: out_word = 8'hFF;
		16'h4940: out_word = 8'hFF;
		16'h4941: out_word = 8'hFF;
		16'h4942: out_word = 8'hFF;
		16'h4943: out_word = 8'hFF;
		16'h4944: out_word = 8'hFF;
		16'h4945: out_word = 8'hFF;
		16'h4946: out_word = 8'hFF;
		16'h4947: out_word = 8'hFF;
		16'h4948: out_word = 8'hFF;
		16'h4949: out_word = 8'hFF;
		16'h494A: out_word = 8'hFF;
		16'h494B: out_word = 8'hFF;
		16'h494C: out_word = 8'hFF;
		16'h494D: out_word = 8'hFF;
		16'h494E: out_word = 8'hFF;
		16'h494F: out_word = 8'hFF;
		16'h4950: out_word = 8'hFF;
		16'h4951: out_word = 8'hFF;
		16'h4952: out_word = 8'hFF;
		16'h4953: out_word = 8'hFF;
		16'h4954: out_word = 8'hFF;
		16'h4955: out_word = 8'hFF;
		16'h4956: out_word = 8'hFF;
		16'h4957: out_word = 8'hFF;
		16'h4958: out_word = 8'hFF;
		16'h4959: out_word = 8'hFF;
		16'h495A: out_word = 8'hFF;
		16'h495B: out_word = 8'hFF;
		16'h495C: out_word = 8'hFF;
		16'h495D: out_word = 8'hFF;
		16'h495E: out_word = 8'hFF;
		16'h495F: out_word = 8'hFF;
		16'h4960: out_word = 8'hFF;
		16'h4961: out_word = 8'hFF;
		16'h4962: out_word = 8'hFF;
		16'h4963: out_word = 8'hFF;
		16'h4964: out_word = 8'hFF;
		16'h4965: out_word = 8'hFF;
		16'h4966: out_word = 8'hFF;
		16'h4967: out_word = 8'hFF;
		16'h4968: out_word = 8'hFF;
		16'h4969: out_word = 8'hFF;
		16'h496A: out_word = 8'hFF;
		16'h496B: out_word = 8'hFF;
		16'h496C: out_word = 8'hFF;
		16'h496D: out_word = 8'hFF;
		16'h496E: out_word = 8'hFF;
		16'h496F: out_word = 8'hFF;
		16'h4970: out_word = 8'hFF;
		16'h4971: out_word = 8'hFF;
		16'h4972: out_word = 8'hFF;
		16'h4973: out_word = 8'hFF;
		16'h4974: out_word = 8'hFF;
		16'h4975: out_word = 8'hFF;
		16'h4976: out_word = 8'hFF;
		16'h4977: out_word = 8'hFF;
		16'h4978: out_word = 8'hFF;
		16'h4979: out_word = 8'hFF;
		16'h497A: out_word = 8'hFF;
		16'h497B: out_word = 8'hFF;
		16'h497C: out_word = 8'hFF;
		16'h497D: out_word = 8'hFF;
		16'h497E: out_word = 8'hFF;
		16'h497F: out_word = 8'hFF;
		16'h4980: out_word = 8'hFF;
		16'h4981: out_word = 8'hFF;
		16'h4982: out_word = 8'hFF;
		16'h4983: out_word = 8'hFF;
		16'h4984: out_word = 8'hFF;
		16'h4985: out_word = 8'hFF;
		16'h4986: out_word = 8'hFF;
		16'h4987: out_word = 8'hFF;
		16'h4988: out_word = 8'hFF;
		16'h4989: out_word = 8'hFF;
		16'h498A: out_word = 8'hFF;
		16'h498B: out_word = 8'hFF;
		16'h498C: out_word = 8'hFF;
		16'h498D: out_word = 8'hFF;
		16'h498E: out_word = 8'hFF;
		16'h498F: out_word = 8'hFF;
		16'h4990: out_word = 8'hFF;
		16'h4991: out_word = 8'hFF;
		16'h4992: out_word = 8'hFF;
		16'h4993: out_word = 8'hFF;
		16'h4994: out_word = 8'hFF;
		16'h4995: out_word = 8'hFF;
		16'h4996: out_word = 8'hFF;
		16'h4997: out_word = 8'hFF;
		16'h4998: out_word = 8'hFF;
		16'h4999: out_word = 8'hFF;
		16'h499A: out_word = 8'hFF;
		16'h499B: out_word = 8'hFF;
		16'h499C: out_word = 8'hFF;
		16'h499D: out_word = 8'hFF;
		16'h499E: out_word = 8'hFF;
		16'h499F: out_word = 8'hFF;
		16'h49A0: out_word = 8'hFF;
		16'h49A1: out_word = 8'hFF;
		16'h49A2: out_word = 8'hFF;
		16'h49A3: out_word = 8'hFF;
		16'h49A4: out_word = 8'hFF;
		16'h49A5: out_word = 8'hFF;
		16'h49A6: out_word = 8'hFF;
		16'h49A7: out_word = 8'hFF;
		16'h49A8: out_word = 8'hFF;
		16'h49A9: out_word = 8'hFF;
		16'h49AA: out_word = 8'hFF;
		16'h49AB: out_word = 8'hFF;
		16'h49AC: out_word = 8'hFF;
		16'h49AD: out_word = 8'hFF;
		16'h49AE: out_word = 8'hFF;
		16'h49AF: out_word = 8'hFF;
		16'h49B0: out_word = 8'hFF;
		16'h49B1: out_word = 8'hFF;
		16'h49B2: out_word = 8'hFF;
		16'h49B3: out_word = 8'hFF;
		16'h49B4: out_word = 8'hFF;
		16'h49B5: out_word = 8'hFF;
		16'h49B6: out_word = 8'hFF;
		16'h49B7: out_word = 8'hFF;
		16'h49B8: out_word = 8'hFF;
		16'h49B9: out_word = 8'hFF;
		16'h49BA: out_word = 8'hFF;
		16'h49BB: out_word = 8'hFF;
		16'h49BC: out_word = 8'hFF;
		16'h49BD: out_word = 8'hFF;
		16'h49BE: out_word = 8'hFF;
		16'h49BF: out_word = 8'hFF;
		16'h49C0: out_word = 8'hFF;
		16'h49C1: out_word = 8'hFF;
		16'h49C2: out_word = 8'hFF;
		16'h49C3: out_word = 8'hFF;
		16'h49C4: out_word = 8'hFF;
		16'h49C5: out_word = 8'hFF;
		16'h49C6: out_word = 8'hFF;
		16'h49C7: out_word = 8'hFF;
		16'h49C8: out_word = 8'hFF;
		16'h49C9: out_word = 8'hFF;
		16'h49CA: out_word = 8'hFF;
		16'h49CB: out_word = 8'hFF;
		16'h49CC: out_word = 8'hFF;
		16'h49CD: out_word = 8'hFF;
		16'h49CE: out_word = 8'hFF;
		16'h49CF: out_word = 8'hFF;
		16'h49D0: out_word = 8'hFF;
		16'h49D1: out_word = 8'hFF;
		16'h49D2: out_word = 8'hFF;
		16'h49D3: out_word = 8'hFF;
		16'h49D4: out_word = 8'hFF;
		16'h49D5: out_word = 8'hFF;
		16'h49D6: out_word = 8'hFF;
		16'h49D7: out_word = 8'hFF;
		16'h49D8: out_word = 8'hFF;
		16'h49D9: out_word = 8'hFF;
		16'h49DA: out_word = 8'hFF;
		16'h49DB: out_word = 8'hFF;
		16'h49DC: out_word = 8'hFF;
		16'h49DD: out_word = 8'hFF;
		16'h49DE: out_word = 8'hFF;
		16'h49DF: out_word = 8'hFF;
		16'h49E0: out_word = 8'hFF;
		16'h49E1: out_word = 8'hFF;
		16'h49E2: out_word = 8'hFF;
		16'h49E3: out_word = 8'hFF;
		16'h49E4: out_word = 8'hFF;
		16'h49E5: out_word = 8'hFF;
		16'h49E6: out_word = 8'hFF;
		16'h49E7: out_word = 8'hFF;
		16'h49E8: out_word = 8'hFF;
		16'h49E9: out_word = 8'hFF;
		16'h49EA: out_word = 8'hFF;
		16'h49EB: out_word = 8'hFF;
		16'h49EC: out_word = 8'hFF;
		16'h49ED: out_word = 8'hFF;
		16'h49EE: out_word = 8'hFF;
		16'h49EF: out_word = 8'hFF;
		16'h49F0: out_word = 8'hFF;
		16'h49F1: out_word = 8'hFF;
		16'h49F2: out_word = 8'hFF;
		16'h49F3: out_word = 8'hFF;
		16'h49F4: out_word = 8'hFF;
		16'h49F5: out_word = 8'hFF;
		16'h49F6: out_word = 8'hFF;
		16'h49F7: out_word = 8'hFF;
		16'h49F8: out_word = 8'hFF;
		16'h49F9: out_word = 8'hFF;
		16'h49FA: out_word = 8'hFF;
		16'h49FB: out_word = 8'hFF;
		16'h49FC: out_word = 8'hFF;
		16'h49FD: out_word = 8'hFF;
		16'h49FE: out_word = 8'hFF;
		16'h49FF: out_word = 8'hFF;
		16'h4A00: out_word = 8'hFF;
		16'h4A01: out_word = 8'h3E;
		16'h4A02: out_word = 8'h3C;
		16'h4A03: out_word = 8'hD3;
		16'h4A04: out_word = 8'hFF;
		16'h4A05: out_word = 8'h3E;
		16'h4A06: out_word = 8'hD0;
		16'h4A07: out_word = 8'hD3;
		16'h4A08: out_word = 8'h1F;
		16'h4A09: out_word = 8'hC9;
		16'h4A0A: out_word = 8'h32;
		16'h4A0B: out_word = 8'h01;
		16'h4A0C: out_word = 8'h5C;
		16'h4A0D: out_word = 8'hF1;
		16'h4A0E: out_word = 8'hC3;
		16'h4A0F: out_word = 8'hC2;
		16'h4A10: out_word = 8'h2E;
		16'h4A11: out_word = 8'h3A;
		16'h4A12: out_word = 8'h01;
		16'h4A13: out_word = 8'h5C;
		16'h4A14: out_word = 8'hED;
		16'h4A15: out_word = 8'h4F;
		16'h4A16: out_word = 8'hF1;
		16'h4A17: out_word = 8'hC3;
		16'h4A18: out_word = 8'h00;
		16'h4A19: out_word = 8'h5C;
		16'h4A1A: out_word = 8'hF5;
		16'h4A1B: out_word = 8'hED;
		16'h4A1C: out_word = 8'h5F;
		16'h4A1D: out_word = 8'hCB;
		16'h4A1E: out_word = 8'h7F;
		16'h4A1F: out_word = 8'h28;
		16'h4A20: out_word = 8'h06;
		16'h4A21: out_word = 8'hD6;
		16'h4A22: out_word = 8'h1F;
		16'h4A23: out_word = 8'hCB;
		16'h4A24: out_word = 8'hFF;
		16'h4A25: out_word = 8'h18;
		16'h4A26: out_word = 8'h04;
		16'h4A27: out_word = 8'hD6;
		16'h4A28: out_word = 8'h1F;
		16'h4A29: out_word = 8'hCB;
		16'h4A2A: out_word = 8'hBF;
		16'h4A2B: out_word = 8'hF5;
		16'h4A2C: out_word = 8'h00;
		16'h4A2D: out_word = 8'h00;
		16'h4A2E: out_word = 8'h00;
		16'h4A2F: out_word = 8'h00;
		16'h4A30: out_word = 8'h00;
		16'h4A31: out_word = 8'h00;
		16'h4A32: out_word = 8'h00;
		16'h4A33: out_word = 8'h00;
		16'h4A34: out_word = 8'h00;
		16'h4A35: out_word = 8'h00;
		16'h4A36: out_word = 8'h00;
		16'h4A37: out_word = 8'h00;
		16'h4A38: out_word = 8'h00;
		16'h4A39: out_word = 8'h00;
		16'h4A3A: out_word = 8'h00;
		16'h4A3B: out_word = 8'h00;
		16'h4A3C: out_word = 8'h00;
		16'h4A3D: out_word = 8'h00;
		16'h4A3E: out_word = 8'h00;
		16'h4A3F: out_word = 8'h00;
		16'h4A40: out_word = 8'h00;
		16'h4A41: out_word = 8'h00;
		16'h4A42: out_word = 8'h00;
		16'h4A43: out_word = 8'h00;
		16'h4A44: out_word = 8'h00;
		16'h4A45: out_word = 8'h3E;
		16'h4A46: out_word = 8'hF7;
		16'h4A47: out_word = 8'hDB;
		16'h4A48: out_word = 8'hFE;
		16'h4A49: out_word = 8'h0F;
		16'h4A4A: out_word = 8'h30;
		16'h4A4B: out_word = 8'h1D;
		16'h4A4C: out_word = 8'h0F;
		16'h4A4D: out_word = 8'h30;
		16'h4A4E: out_word = 8'h20;
		16'h4A4F: out_word = 8'h0F;
		16'h4A50: out_word = 8'h30;
		16'h4A51: out_word = 8'h2C;
		16'h4A52: out_word = 8'h0F;
		16'h4A53: out_word = 8'h38;
		16'h4A54: out_word = 8'hF0;
		16'h4A55: out_word = 8'hF1;
		16'h4A56: out_word = 8'hCB;
		16'h4A57: out_word = 8'h7F;
		16'h4A58: out_word = 8'h28;
		16'h4A59: out_word = 8'h06;
		16'h4A5A: out_word = 8'hC6;
		16'h4A5B: out_word = 8'h17;
		16'h4A5C: out_word = 8'hCB;
		16'h4A5D: out_word = 8'hFF;
		16'h4A5E: out_word = 8'h18;
		16'h4A5F: out_word = 8'h04;
		16'h4A60: out_word = 8'hC6;
		16'h4A61: out_word = 8'h17;
		16'h4A62: out_word = 8'hCB;
		16'h4A63: out_word = 8'hBF;
		16'h4A64: out_word = 8'hED;
		16'h4A65: out_word = 8'h4F;
		16'h4A66: out_word = 8'hF1;
		16'h4A67: out_word = 8'hED;
		16'h4A68: out_word = 8'h45;
		16'h4A69: out_word = 8'hF1;
		16'h4A6A: out_word = 8'hED;
		16'h4A6B: out_word = 8'h4F;
		16'h4A6C: out_word = 8'hF1;
		16'h4A6D: out_word = 8'h18;
		16'h4A6E: out_word = 8'h09;
		16'h4A6F: out_word = 8'hF1;
		16'h4A70: out_word = 8'hF1;
		16'h4A71: out_word = 8'hED;
		16'h4A72: out_word = 8'h73;
		16'h4A73: out_word = 8'hFE;
		16'h4A74: out_word = 8'h57;
		16'h4A75: out_word = 8'h31;
		16'h4A76: out_word = 8'h00;
		16'h4A77: out_word = 8'h58;
		16'h4A78: out_word = 8'hF5;
		16'h4A79: out_word = 8'hC5;
		16'h4A7A: out_word = 8'hD5;
		16'h4A7B: out_word = 8'hC3;
		16'h4A7C: out_word = 8'h59;
		16'h4A7D: out_word = 8'h2A;
		16'h4A7E: out_word = 8'hF1;
		16'h4A7F: out_word = 8'hED;
		16'h4A80: out_word = 8'h4F;
		16'h4A81: out_word = 8'hE5;
		16'h4A82: out_word = 8'h21;
		16'h4A83: out_word = 8'h00;
		16'h4A84: out_word = 8'h00;
		16'h4A85: out_word = 8'h39;
		16'h4A86: out_word = 8'h23;
		16'h4A87: out_word = 8'h23;
		16'h4A88: out_word = 8'h7C;
		16'h4A89: out_word = 8'hE1;
		16'h4A8A: out_word = 8'hFE;
		16'h4A8B: out_word = 8'hC0;
		16'h4A8C: out_word = 8'h30;
		16'h4A8D: out_word = 8'h36;
		16'h4A8E: out_word = 8'hED;
		16'h4A8F: out_word = 8'h5F;
		16'h4A90: out_word = 8'hCB;
		16'h4A91: out_word = 8'h7F;
		16'h4A92: out_word = 8'h28;
		16'h4A93: out_word = 8'h06;
		16'h4A94: out_word = 8'hD6;
		16'h4A95: out_word = 8'h09;
		16'h4A96: out_word = 8'hCB;
		16'h4A97: out_word = 8'hFF;
		16'h4A98: out_word = 8'h18;
		16'h4A99: out_word = 8'h04;
		16'h4A9A: out_word = 8'hD6;
		16'h4A9B: out_word = 8'h09;
		16'h4A9C: out_word = 8'hCB;
		16'h4A9D: out_word = 8'hBF;
		16'h4A9E: out_word = 8'hED;
		16'h4A9F: out_word = 8'h4F;
		16'h4AA0: out_word = 8'hC5;
		16'h4AA1: out_word = 8'h01;
		16'h4AA2: out_word = 8'hFD;
		16'h4AA3: out_word = 8'hFF;
		16'h4AA4: out_word = 8'h3E;
		16'h4AA5: out_word = 8'h07;
		16'h4AA6: out_word = 8'hED;
		16'h4AA7: out_word = 8'h79;
		16'h4AA8: out_word = 8'h06;
		16'h4AA9: out_word = 8'hBF;
		16'h4AAA: out_word = 8'h3E;
		16'h4AAB: out_word = 8'hFF;
		16'h4AAC: out_word = 8'hED;
		16'h4AAD: out_word = 8'h79;
		16'h4AAE: out_word = 8'h3E;
		16'h4AAF: out_word = 8'h57;
		16'h4AB0: out_word = 8'h01;
		16'h4AB1: out_word = 8'hFD;
		16'h4AB2: out_word = 8'h7F;
		16'h4AB3: out_word = 8'hED;
		16'h4AB4: out_word = 8'h79;
		16'h4AB5: out_word = 8'hC1;
		16'h4AB6: out_word = 8'hF1;
		16'h4AB7: out_word = 8'hE3;
		16'h4AB8: out_word = 8'h22;
		16'h4AB9: out_word = 8'hE4;
		16'h4ABA: out_word = 8'hFE;
		16'h4ABB: out_word = 8'h22;
		16'h4ABC: out_word = 8'hFE;
		16'h4ABD: out_word = 8'hFE;
		16'h4ABE: out_word = 8'hE3;
		16'h4ABF: out_word = 8'h33;
		16'h4AC0: out_word = 8'h33;
		16'h4AC1: out_word = 8'hC3;
		16'h4AC2: out_word = 8'h00;
		16'h4AC3: out_word = 8'hDB;
		16'h4AC4: out_word = 8'hED;
		16'h4AC5: out_word = 8'h5F;
		16'h4AC6: out_word = 8'hCB;
		16'h4AC7: out_word = 8'h7F;
		16'h4AC8: out_word = 8'h28;
		16'h4AC9: out_word = 8'h06;
		16'h4ACA: out_word = 8'hD6;
		16'h4ACB: out_word = 8'h15;
		16'h4ACC: out_word = 8'hCB;
		16'h4ACD: out_word = 8'hFF;
		16'h4ACE: out_word = 8'h18;
		16'h4ACF: out_word = 8'h04;
		16'h4AD0: out_word = 8'hD6;
		16'h4AD1: out_word = 8'h15;
		16'h4AD2: out_word = 8'hCB;
		16'h4AD3: out_word = 8'hBF;
		16'h4AD4: out_word = 8'hED;
		16'h4AD5: out_word = 8'h4F;
		16'h4AD6: out_word = 8'hF1;
		16'h4AD7: out_word = 8'hED;
		16'h4AD8: out_word = 8'h73;
		16'h4AD9: out_word = 8'h00;
		16'h4ADA: out_word = 8'h58;
		16'h4ADB: out_word = 8'hE3;
		16'h4ADC: out_word = 8'h22;
		16'h4ADD: out_word = 8'h02;
		16'h4ADE: out_word = 8'h58;
		16'h4ADF: out_word = 8'hE3;
		16'h4AE0: out_word = 8'h31;
		16'h4AE1: out_word = 8'h08;
		16'h4AE2: out_word = 8'h58;
		16'h4AE3: out_word = 8'hF5;
		16'h4AE4: out_word = 8'hC5;
		16'h4AE5: out_word = 8'h01;
		16'h4AE6: out_word = 8'hFD;
		16'h4AE7: out_word = 8'hFF;
		16'h4AE8: out_word = 8'h3E;
		16'h4AE9: out_word = 8'h07;
		16'h4AEA: out_word = 8'hED;
		16'h4AEB: out_word = 8'h79;
		16'h4AEC: out_word = 8'h06;
		16'h4AED: out_word = 8'hBF;
		16'h4AEE: out_word = 8'h3E;
		16'h4AEF: out_word = 8'hFF;
		16'h4AF0: out_word = 8'hED;
		16'h4AF1: out_word = 8'h79;
		16'h4AF2: out_word = 8'h3E;
		16'h4AF3: out_word = 8'h57;
		16'h4AF4: out_word = 8'h01;
		16'h4AF5: out_word = 8'hFD;
		16'h4AF6: out_word = 8'h7F;
		16'h4AF7: out_word = 8'hED;
		16'h4AF8: out_word = 8'h79;
		16'h4AF9: out_word = 8'hC1;
		16'h4AFA: out_word = 8'hF1;
		16'h4AFB: out_word = 8'hED;
		16'h4AFC: out_word = 8'h7B;
		16'h4AFD: out_word = 8'h00;
		16'h4AFE: out_word = 8'h58;
		16'h4AFF: out_word = 8'h22;
		16'h4B00: out_word = 8'h00;
		16'h4B01: out_word = 8'hC0;
		16'h4B02: out_word = 8'h2A;
		16'h4B03: out_word = 8'h02;
		16'h4B04: out_word = 8'h58;
		16'h4B05: out_word = 8'h22;
		16'h4B06: out_word = 8'hE4;
		16'h4B07: out_word = 8'hFE;
		16'h4B08: out_word = 8'h22;
		16'h4B09: out_word = 8'hFE;
		16'h4B0A: out_word = 8'hFE;
		16'h4B0B: out_word = 8'h2A;
		16'h4B0C: out_word = 8'h00;
		16'h4B0D: out_word = 8'hC0;
		16'h4B0E: out_word = 8'h18;
		16'h4B0F: out_word = 8'hAF;
		16'h4B10: out_word = 8'hFF;
		16'h4B11: out_word = 8'hFF;
		16'h4B12: out_word = 8'hFF;
		16'h4B13: out_word = 8'hFF;
		16'h4B14: out_word = 8'hFF;
		16'h4B15: out_word = 8'hFF;
		16'h4B16: out_word = 8'hFF;
		16'h4B17: out_word = 8'hFF;
		16'h4B18: out_word = 8'hFF;
		16'h4B19: out_word = 8'hFF;
		16'h4B1A: out_word = 8'hFF;
		16'h4B1B: out_word = 8'hFF;
		16'h4B1C: out_word = 8'hFF;
		16'h4B1D: out_word = 8'hFF;
		16'h4B1E: out_word = 8'hFF;
		16'h4B1F: out_word = 8'hFF;
		16'h4B20: out_word = 8'hFF;
		16'h4B21: out_word = 8'hFF;
		16'h4B22: out_word = 8'hFF;
		16'h4B23: out_word = 8'hFF;
		16'h4B24: out_word = 8'hFF;
		16'h4B25: out_word = 8'hFF;
		16'h4B26: out_word = 8'hFF;
		16'h4B27: out_word = 8'hFF;
		16'h4B28: out_word = 8'hFF;
		16'h4B29: out_word = 8'hFF;
		16'h4B2A: out_word = 8'hFF;
		16'h4B2B: out_word = 8'hFF;
		16'h4B2C: out_word = 8'hFF;
		16'h4B2D: out_word = 8'hFF;
		16'h4B2E: out_word = 8'hFF;
		16'h4B2F: out_word = 8'hFF;
		16'h4B30: out_word = 8'hFF;
		16'h4B31: out_word = 8'hFF;
		16'h4B32: out_word = 8'hFF;
		16'h4B33: out_word = 8'hFF;
		16'h4B34: out_word = 8'hFF;
		16'h4B35: out_word = 8'hFF;
		16'h4B36: out_word = 8'hFF;
		16'h4B37: out_word = 8'hFF;
		16'h4B38: out_word = 8'hFF;
		16'h4B39: out_word = 8'hFF;
		16'h4B3A: out_word = 8'hFF;
		16'h4B3B: out_word = 8'hFF;
		16'h4B3C: out_word = 8'hFF;
		16'h4B3D: out_word = 8'hFF;
		16'h4B3E: out_word = 8'hFF;
		16'h4B3F: out_word = 8'hFF;
		16'h4B40: out_word = 8'hFF;
		16'h4B41: out_word = 8'hFF;
		16'h4B42: out_word = 8'hFF;
		16'h4B43: out_word = 8'hFF;
		16'h4B44: out_word = 8'hFF;
		16'h4B45: out_word = 8'hFF;
		16'h4B46: out_word = 8'hFF;
		16'h4B47: out_word = 8'hFF;
		16'h4B48: out_word = 8'hFF;
		16'h4B49: out_word = 8'hFF;
		16'h4B4A: out_word = 8'hFF;
		16'h4B4B: out_word = 8'hFF;
		16'h4B4C: out_word = 8'hFF;
		16'h4B4D: out_word = 8'hFF;
		16'h4B4E: out_word = 8'hFF;
		16'h4B4F: out_word = 8'hFF;
		16'h4B50: out_word = 8'hFF;
		16'h4B51: out_word = 8'hFF;
		16'h4B52: out_word = 8'hFF;
		16'h4B53: out_word = 8'hFF;
		16'h4B54: out_word = 8'hFF;
		16'h4B55: out_word = 8'hFF;
		16'h4B56: out_word = 8'hFF;
		16'h4B57: out_word = 8'hFF;
		16'h4B58: out_word = 8'hFF;
		16'h4B59: out_word = 8'hFF;
		16'h4B5A: out_word = 8'hFF;
		16'h4B5B: out_word = 8'hFF;
		16'h4B5C: out_word = 8'hFF;
		16'h4B5D: out_word = 8'hFF;
		16'h4B5E: out_word = 8'hFF;
		16'h4B5F: out_word = 8'hFF;
		16'h4B60: out_word = 8'hFF;
		16'h4B61: out_word = 8'hFF;
		16'h4B62: out_word = 8'hFF;
		16'h4B63: out_word = 8'hFF;
		16'h4B64: out_word = 8'hFF;
		16'h4B65: out_word = 8'hFF;
		16'h4B66: out_word = 8'hFF;
		16'h4B67: out_word = 8'hFF;
		16'h4B68: out_word = 8'hFF;
		16'h4B69: out_word = 8'hFF;
		16'h4B6A: out_word = 8'hFF;
		16'h4B6B: out_word = 8'hFF;
		16'h4B6C: out_word = 8'hFF;
		16'h4B6D: out_word = 8'hFF;
		16'h4B6E: out_word = 8'hFF;
		16'h4B6F: out_word = 8'hFF;
		16'h4B70: out_word = 8'hFF;
		16'h4B71: out_word = 8'hFF;
		16'h4B72: out_word = 8'hFF;
		16'h4B73: out_word = 8'hFF;
		16'h4B74: out_word = 8'hFF;
		16'h4B75: out_word = 8'hFF;
		16'h4B76: out_word = 8'hFF;
		16'h4B77: out_word = 8'hFF;
		16'h4B78: out_word = 8'hFF;
		16'h4B79: out_word = 8'hFF;
		16'h4B7A: out_word = 8'hFF;
		16'h4B7B: out_word = 8'hFF;
		16'h4B7C: out_word = 8'hFF;
		16'h4B7D: out_word = 8'hFF;
		16'h4B7E: out_word = 8'hFF;
		16'h4B7F: out_word = 8'hFF;
		16'h4B80: out_word = 8'hFF;
		16'h4B81: out_word = 8'hFF;
		16'h4B82: out_word = 8'hFF;
		16'h4B83: out_word = 8'hFF;
		16'h4B84: out_word = 8'hFF;
		16'h4B85: out_word = 8'hFF;
		16'h4B86: out_word = 8'hFF;
		16'h4B87: out_word = 8'hFF;
		16'h4B88: out_word = 8'hFF;
		16'h4B89: out_word = 8'hFF;
		16'h4B8A: out_word = 8'hFF;
		16'h4B8B: out_word = 8'hFF;
		16'h4B8C: out_word = 8'hFF;
		16'h4B8D: out_word = 8'hFF;
		16'h4B8E: out_word = 8'hFF;
		16'h4B8F: out_word = 8'hFF;
		16'h4B90: out_word = 8'hFF;
		16'h4B91: out_word = 8'hFF;
		16'h4B92: out_word = 8'hFF;
		16'h4B93: out_word = 8'hFF;
		16'h4B94: out_word = 8'hFF;
		16'h4B95: out_word = 8'hFF;
		16'h4B96: out_word = 8'hFF;
		16'h4B97: out_word = 8'hFF;
		16'h4B98: out_word = 8'hFF;
		16'h4B99: out_word = 8'hFF;
		16'h4B9A: out_word = 8'hFF;
		16'h4B9B: out_word = 8'hFF;
		16'h4B9C: out_word = 8'hFF;
		16'h4B9D: out_word = 8'hFF;
		16'h4B9E: out_word = 8'hFF;
		16'h4B9F: out_word = 8'hFF;
		16'h4BA0: out_word = 8'hFF;
		16'h4BA1: out_word = 8'hFF;
		16'h4BA2: out_word = 8'hFF;
		16'h4BA3: out_word = 8'hFF;
		16'h4BA4: out_word = 8'hFF;
		16'h4BA5: out_word = 8'hFF;
		16'h4BA6: out_word = 8'hFF;
		16'h4BA7: out_word = 8'hFF;
		16'h4BA8: out_word = 8'hFF;
		16'h4BA9: out_word = 8'hFF;
		16'h4BAA: out_word = 8'hFF;
		16'h4BAB: out_word = 8'hFF;
		16'h4BAC: out_word = 8'hFF;
		16'h4BAD: out_word = 8'hFF;
		16'h4BAE: out_word = 8'hFF;
		16'h4BAF: out_word = 8'hFF;
		16'h4BB0: out_word = 8'hFF;
		16'h4BB1: out_word = 8'hFF;
		16'h4BB2: out_word = 8'hFF;
		16'h4BB3: out_word = 8'hFF;
		16'h4BB4: out_word = 8'hFF;
		16'h4BB5: out_word = 8'hFF;
		16'h4BB6: out_word = 8'hFF;
		16'h4BB7: out_word = 8'hFF;
		16'h4BB8: out_word = 8'hFF;
		16'h4BB9: out_word = 8'hFF;
		16'h4BBA: out_word = 8'hFF;
		16'h4BBB: out_word = 8'hFF;
		16'h4BBC: out_word = 8'hFF;
		16'h4BBD: out_word = 8'hFF;
		16'h4BBE: out_word = 8'hFF;
		16'h4BBF: out_word = 8'hFF;
		16'h4BC0: out_word = 8'hFF;
		16'h4BC1: out_word = 8'hFF;
		16'h4BC2: out_word = 8'hFF;
		16'h4BC3: out_word = 8'hFF;
		16'h4BC4: out_word = 8'hFF;
		16'h4BC5: out_word = 8'hFF;
		16'h4BC6: out_word = 8'hFF;
		16'h4BC7: out_word = 8'hFF;
		16'h4BC8: out_word = 8'hFF;
		16'h4BC9: out_word = 8'hFF;
		16'h4BCA: out_word = 8'hFF;
		16'h4BCB: out_word = 8'hFF;
		16'h4BCC: out_word = 8'hFF;
		16'h4BCD: out_word = 8'hFF;
		16'h4BCE: out_word = 8'hFF;
		16'h4BCF: out_word = 8'hFF;
		16'h4BD0: out_word = 8'hFF;
		16'h4BD1: out_word = 8'hFF;
		16'h4BD2: out_word = 8'hFF;
		16'h4BD3: out_word = 8'hFF;
		16'h4BD4: out_word = 8'hFF;
		16'h4BD5: out_word = 8'hFF;
		16'h4BD6: out_word = 8'hFF;
		16'h4BD7: out_word = 8'hFF;
		16'h4BD8: out_word = 8'hFF;
		16'h4BD9: out_word = 8'hFF;
		16'h4BDA: out_word = 8'hFF;
		16'h4BDB: out_word = 8'hFF;
		16'h4BDC: out_word = 8'hFF;
		16'h4BDD: out_word = 8'hFF;
		16'h4BDE: out_word = 8'hFF;
		16'h4BDF: out_word = 8'hFF;
		16'h4BE0: out_word = 8'hFF;
		16'h4BE1: out_word = 8'hFF;
		16'h4BE2: out_word = 8'hFF;
		16'h4BE3: out_word = 8'hFF;
		16'h4BE4: out_word = 8'hFF;
		16'h4BE5: out_word = 8'hFF;
		16'h4BE6: out_word = 8'hFF;
		16'h4BE7: out_word = 8'hFF;
		16'h4BE8: out_word = 8'hFF;
		16'h4BE9: out_word = 8'hFF;
		16'h4BEA: out_word = 8'hFF;
		16'h4BEB: out_word = 8'hFF;
		16'h4BEC: out_word = 8'hFF;
		16'h4BED: out_word = 8'hFF;
		16'h4BEE: out_word = 8'hFF;
		16'h4BEF: out_word = 8'hFF;
		16'h4BF0: out_word = 8'hFF;
		16'h4BF1: out_word = 8'hFF;
		16'h4BF2: out_word = 8'hFF;
		16'h4BF3: out_word = 8'hFF;
		16'h4BF4: out_word = 8'hFF;
		16'h4BF5: out_word = 8'hFF;
		16'h4BF6: out_word = 8'hFF;
		16'h4BF7: out_word = 8'hFF;
		16'h4BF8: out_word = 8'hFF;
		16'h4BF9: out_word = 8'hFF;
		16'h4BFA: out_word = 8'hFF;
		16'h4BFB: out_word = 8'hFF;
		16'h4BFC: out_word = 8'hFF;
		16'h4BFD: out_word = 8'hFF;
		16'h4BFE: out_word = 8'hFF;
		16'h4BFF: out_word = 8'hFF;
		16'h4C00: out_word = 8'h00;
		16'h4C01: out_word = 8'h00;
		16'h4C02: out_word = 8'h4C;
		16'h4C03: out_word = 8'h52;
		16'h4C04: out_word = 8'h72;
		16'h4C05: out_word = 8'h52;
		16'h4C06: out_word = 8'h4C;
		16'h4C07: out_word = 8'h00;
		16'h4C08: out_word = 8'h00;
		16'h4C09: out_word = 8'h00;
		16'h4C0A: out_word = 8'h38;
		16'h4C0B: out_word = 8'h04;
		16'h4C0C: out_word = 8'h3C;
		16'h4C0D: out_word = 8'h44;
		16'h4C0E: out_word = 8'h3C;
		16'h4C0F: out_word = 8'h00;
		16'h4C10: out_word = 8'h00;
		16'h4C11: out_word = 8'h00;
		16'h4C12: out_word = 8'h78;
		16'h4C13: out_word = 8'h40;
		16'h4C14: out_word = 8'h78;
		16'h4C15: out_word = 8'h44;
		16'h4C16: out_word = 8'h78;
		16'h4C17: out_word = 8'h00;
		16'h4C18: out_word = 8'h00;
		16'h4C19: out_word = 8'h00;
		16'h4C1A: out_word = 8'h48;
		16'h4C1B: out_word = 8'h48;
		16'h4C1C: out_word = 8'h48;
		16'h4C1D: out_word = 8'h48;
		16'h4C1E: out_word = 8'h7C;
		16'h4C1F: out_word = 8'h04;
		16'h4C20: out_word = 8'h00;
		16'h4C21: out_word = 8'h00;
		16'h4C22: out_word = 8'h18;
		16'h4C23: out_word = 8'h28;
		16'h4C24: out_word = 8'h28;
		16'h4C25: out_word = 8'h28;
		16'h4C26: out_word = 8'h7C;
		16'h4C27: out_word = 8'h44;
		16'h4C28: out_word = 8'h00;
		16'h4C29: out_word = 8'h00;
		16'h4C2A: out_word = 8'h38;
		16'h4C2B: out_word = 8'h44;
		16'h4C2C: out_word = 8'h78;
		16'h4C2D: out_word = 8'h40;
		16'h4C2E: out_word = 8'h3C;
		16'h4C2F: out_word = 8'h00;
		16'h4C30: out_word = 8'h00;
		16'h4C31: out_word = 8'h10;
		16'h4C32: out_word = 8'h38;
		16'h4C33: out_word = 8'h54;
		16'h4C34: out_word = 8'h54;
		16'h4C35: out_word = 8'h38;
		16'h4C36: out_word = 8'h10;
		16'h4C37: out_word = 8'h00;
		16'h4C38: out_word = 8'h00;
		16'h4C39: out_word = 8'h00;
		16'h4C3A: out_word = 8'h7C;
		16'h4C3B: out_word = 8'h40;
		16'h4C3C: out_word = 8'h40;
		16'h4C3D: out_word = 8'h40;
		16'h4C3E: out_word = 8'h40;
		16'h4C3F: out_word = 8'h00;
		16'h4C40: out_word = 8'h00;
		16'h4C41: out_word = 8'h00;
		16'h4C42: out_word = 8'h44;
		16'h4C43: out_word = 8'h28;
		16'h4C44: out_word = 8'h10;
		16'h4C45: out_word = 8'h28;
		16'h4C46: out_word = 8'h44;
		16'h4C47: out_word = 8'h00;
		16'h4C48: out_word = 8'h00;
		16'h4C49: out_word = 8'h00;
		16'h4C4A: out_word = 8'h44;
		16'h4C4B: out_word = 8'h4C;
		16'h4C4C: out_word = 8'h54;
		16'h4C4D: out_word = 8'h64;
		16'h4C4E: out_word = 8'h44;
		16'h4C4F: out_word = 8'h00;
		16'h4C50: out_word = 8'h00;
		16'h4C51: out_word = 8'h10;
		16'h4C52: out_word = 8'h44;
		16'h4C53: out_word = 8'h4C;
		16'h4C54: out_word = 8'h54;
		16'h4C55: out_word = 8'h64;
		16'h4C56: out_word = 8'h44;
		16'h4C57: out_word = 8'h00;
		16'h4C58: out_word = 8'h00;
		16'h4C59: out_word = 8'h00;
		16'h4C5A: out_word = 8'h48;
		16'h4C5B: out_word = 8'h50;
		16'h4C5C: out_word = 8'h70;
		16'h4C5D: out_word = 8'h48;
		16'h4C5E: out_word = 8'h44;
		16'h4C5F: out_word = 8'h00;
		16'h4C60: out_word = 8'h00;
		16'h4C61: out_word = 8'h00;
		16'h4C62: out_word = 8'h1C;
		16'h4C63: out_word = 8'h24;
		16'h4C64: out_word = 8'h24;
		16'h4C65: out_word = 8'h24;
		16'h4C66: out_word = 8'h44;
		16'h4C67: out_word = 8'h00;
		16'h4C68: out_word = 8'h00;
		16'h4C69: out_word = 8'h00;
		16'h4C6A: out_word = 8'h44;
		16'h4C6B: out_word = 8'h6C;
		16'h4C6C: out_word = 8'h54;
		16'h4C6D: out_word = 8'h54;
		16'h4C6E: out_word = 8'h44;
		16'h4C6F: out_word = 8'h00;
		16'h4C70: out_word = 8'h00;
		16'h4C71: out_word = 8'h00;
		16'h4C72: out_word = 8'h44;
		16'h4C73: out_word = 8'h44;
		16'h4C74: out_word = 8'h7C;
		16'h4C75: out_word = 8'h44;
		16'h4C76: out_word = 8'h44;
		16'h4C77: out_word = 8'h00;
		16'h4C78: out_word = 8'h00;
		16'h4C79: out_word = 8'h00;
		16'h4C7A: out_word = 8'h38;
		16'h4C7B: out_word = 8'h44;
		16'h4C7C: out_word = 8'h44;
		16'h4C7D: out_word = 8'h44;
		16'h4C7E: out_word = 8'h38;
		16'h4C7F: out_word = 8'h00;
		16'h4C80: out_word = 8'h00;
		16'h4C81: out_word = 8'h00;
		16'h4C82: out_word = 8'h7C;
		16'h4C83: out_word = 8'h44;
		16'h4C84: out_word = 8'h44;
		16'h4C85: out_word = 8'h44;
		16'h4C86: out_word = 8'h44;
		16'h4C87: out_word = 8'h00;
		16'h4C88: out_word = 8'h00;
		16'h4C89: out_word = 8'h00;
		16'h4C8A: out_word = 8'h3C;
		16'h4C8B: out_word = 8'h44;
		16'h4C8C: out_word = 8'h3C;
		16'h4C8D: out_word = 8'h24;
		16'h4C8E: out_word = 8'h44;
		16'h4C8F: out_word = 8'h00;
		16'h4C90: out_word = 8'h00;
		16'h4C91: out_word = 8'h00;
		16'h4C92: out_word = 8'h78;
		16'h4C93: out_word = 8'h44;
		16'h4C94: out_word = 8'h44;
		16'h4C95: out_word = 8'h78;
		16'h4C96: out_word = 8'h40;
		16'h4C97: out_word = 8'h40;
		16'h4C98: out_word = 8'h00;
		16'h4C99: out_word = 8'h00;
		16'h4C9A: out_word = 8'h38;
		16'h4C9B: out_word = 8'h40;
		16'h4C9C: out_word = 8'h40;
		16'h4C9D: out_word = 8'h40;
		16'h4C9E: out_word = 8'h38;
		16'h4C9F: out_word = 8'h00;
		16'h4CA0: out_word = 8'h00;
		16'h4CA1: out_word = 8'h00;
		16'h4CA2: out_word = 8'h7C;
		16'h4CA3: out_word = 8'h10;
		16'h4CA4: out_word = 8'h10;
		16'h4CA5: out_word = 8'h10;
		16'h4CA6: out_word = 8'h10;
		16'h4CA7: out_word = 8'h00;
		16'h4CA8: out_word = 8'h00;
		16'h4CA9: out_word = 8'h00;
		16'h4CAA: out_word = 8'h44;
		16'h4CAB: out_word = 8'h44;
		16'h4CAC: out_word = 8'h3C;
		16'h4CAD: out_word = 8'h04;
		16'h4CAE: out_word = 8'h38;
		16'h4CAF: out_word = 8'h00;
		16'h4CB0: out_word = 8'h00;
		16'h4CB1: out_word = 8'h00;
		16'h4CB2: out_word = 8'h54;
		16'h4CB3: out_word = 8'h54;
		16'h4CB4: out_word = 8'h38;
		16'h4CB5: out_word = 8'h54;
		16'h4CB6: out_word = 8'h54;
		16'h4CB7: out_word = 8'h00;
		16'h4CB8: out_word = 8'h00;
		16'h4CB9: out_word = 8'h00;
		16'h4CBA: out_word = 8'h78;
		16'h4CBB: out_word = 8'h44;
		16'h4CBC: out_word = 8'h78;
		16'h4CBD: out_word = 8'h44;
		16'h4CBE: out_word = 8'h78;
		16'h4CBF: out_word = 8'h00;
		16'h4CC0: out_word = 8'h00;
		16'h4CC1: out_word = 8'h00;
		16'h4CC2: out_word = 8'h40;
		16'h4CC3: out_word = 8'h40;
		16'h4CC4: out_word = 8'h78;
		16'h4CC5: out_word = 8'h44;
		16'h4CC6: out_word = 8'h78;
		16'h4CC7: out_word = 8'h00;
		16'h4CC8: out_word = 8'h00;
		16'h4CC9: out_word = 8'h00;
		16'h4CCA: out_word = 8'h44;
		16'h4CCB: out_word = 8'h44;
		16'h4CCC: out_word = 8'h74;
		16'h4CCD: out_word = 8'h4C;
		16'h4CCE: out_word = 8'h74;
		16'h4CCF: out_word = 8'h00;
		16'h4CD0: out_word = 8'h00;
		16'h4CD1: out_word = 8'h00;
		16'h4CD2: out_word = 8'h38;
		16'h4CD3: out_word = 8'h44;
		16'h4CD4: out_word = 8'h18;
		16'h4CD5: out_word = 8'h44;
		16'h4CD6: out_word = 8'h38;
		16'h4CD7: out_word = 8'h00;
		16'h4CD8: out_word = 8'h00;
		16'h4CD9: out_word = 8'h00;
		16'h4CDA: out_word = 8'h54;
		16'h4CDB: out_word = 8'h54;
		16'h4CDC: out_word = 8'h54;
		16'h4CDD: out_word = 8'h54;
		16'h4CDE: out_word = 8'h7C;
		16'h4CDF: out_word = 8'h00;
		16'h4CE0: out_word = 8'h00;
		16'h4CE1: out_word = 8'h00;
		16'h4CE2: out_word = 8'h38;
		16'h4CE3: out_word = 8'h04;
		16'h4CE4: out_word = 8'h1C;
		16'h4CE5: out_word = 8'h04;
		16'h4CE6: out_word = 8'h38;
		16'h4CE7: out_word = 8'h00;
		16'h4CE8: out_word = 8'h00;
		16'h4CE9: out_word = 8'h00;
		16'h4CEA: out_word = 8'h54;
		16'h4CEB: out_word = 8'h54;
		16'h4CEC: out_word = 8'h54;
		16'h4CED: out_word = 8'h54;
		16'h4CEE: out_word = 8'h7E;
		16'h4CEF: out_word = 8'h02;
		16'h4CF0: out_word = 8'h00;
		16'h4CF1: out_word = 8'h00;
		16'h4CF2: out_word = 8'h44;
		16'h4CF3: out_word = 8'h44;
		16'h4CF4: out_word = 8'h3C;
		16'h4CF5: out_word = 8'h04;
		16'h4CF6: out_word = 8'h04;
		16'h4CF7: out_word = 8'h00;
		16'h4CF8: out_word = 8'h00;
		16'h4CF9: out_word = 8'h00;
		16'h4CFA: out_word = 8'h60;
		16'h4CFB: out_word = 8'h20;
		16'h4CFC: out_word = 8'h38;
		16'h4CFD: out_word = 8'h24;
		16'h4CFE: out_word = 8'h38;
		16'h4CFF: out_word = 8'h00;
		16'h4D00: out_word = 8'h00;
		16'h4D01: out_word = 8'h4C;
		16'h4D02: out_word = 8'h52;
		16'h4D03: out_word = 8'h72;
		16'h4D04: out_word = 8'h52;
		16'h4D05: out_word = 8'h52;
		16'h4D06: out_word = 8'h4C;
		16'h4D07: out_word = 8'h00;
		16'h4D08: out_word = 8'h00;
		16'h4D09: out_word = 8'h3C;
		16'h4D0A: out_word = 8'h42;
		16'h4D0B: out_word = 8'h42;
		16'h4D0C: out_word = 8'h7E;
		16'h4D0D: out_word = 8'h42;
		16'h4D0E: out_word = 8'h42;
		16'h4D0F: out_word = 8'h00;
		16'h4D10: out_word = 8'h00;
		16'h4D11: out_word = 8'h7C;
		16'h4D12: out_word = 8'h40;
		16'h4D13: out_word = 8'h7C;
		16'h4D14: out_word = 8'h42;
		16'h4D15: out_word = 8'h42;
		16'h4D16: out_word = 8'h7C;
		16'h4D17: out_word = 8'h00;
		16'h4D18: out_word = 8'h00;
		16'h4D19: out_word = 8'h44;
		16'h4D1A: out_word = 8'h44;
		16'h4D1B: out_word = 8'h44;
		16'h4D1C: out_word = 8'h44;
		16'h4D1D: out_word = 8'h44;
		16'h4D1E: out_word = 8'h7E;
		16'h4D1F: out_word = 8'h02;
		16'h4D20: out_word = 8'h00;
		16'h4D21: out_word = 8'h18;
		16'h4D22: out_word = 8'h24;
		16'h4D23: out_word = 8'h24;
		16'h4D24: out_word = 8'h24;
		16'h4D25: out_word = 8'h24;
		16'h4D26: out_word = 8'h7E;
		16'h4D27: out_word = 8'h42;
		16'h4D28: out_word = 8'h00;
		16'h4D29: out_word = 8'h7E;
		16'h4D2A: out_word = 8'h40;
		16'h4D2B: out_word = 8'h7C;
		16'h4D2C: out_word = 8'h40;
		16'h4D2D: out_word = 8'h40;
		16'h4D2E: out_word = 8'h7E;
		16'h4D2F: out_word = 8'h00;
		16'h4D30: out_word = 8'h00;
		16'h4D31: out_word = 8'h38;
		16'h4D32: out_word = 8'h54;
		16'h4D33: out_word = 8'h54;
		16'h4D34: out_word = 8'h38;
		16'h4D35: out_word = 8'h10;
		16'h4D36: out_word = 8'h10;
		16'h4D37: out_word = 8'h00;
		16'h4D38: out_word = 8'h00;
		16'h4D39: out_word = 8'h7E;
		16'h4D3A: out_word = 8'h40;
		16'h4D3B: out_word = 8'h40;
		16'h4D3C: out_word = 8'h40;
		16'h4D3D: out_word = 8'h40;
		16'h4D3E: out_word = 8'h40;
		16'h4D3F: out_word = 8'h00;
		16'h4D40: out_word = 8'h00;
		16'h4D41: out_word = 8'h42;
		16'h4D42: out_word = 8'h24;
		16'h4D43: out_word = 8'h18;
		16'h4D44: out_word = 8'h18;
		16'h4D45: out_word = 8'h24;
		16'h4D46: out_word = 8'h42;
		16'h4D47: out_word = 8'h00;
		16'h4D48: out_word = 8'h00;
		16'h4D49: out_word = 8'h42;
		16'h4D4A: out_word = 8'h46;
		16'h4D4B: out_word = 8'h4A;
		16'h4D4C: out_word = 8'h52;
		16'h4D4D: out_word = 8'h62;
		16'h4D4E: out_word = 8'h42;
		16'h4D4F: out_word = 8'h00;
		16'h4D50: out_word = 8'h00;
		16'h4D51: out_word = 8'h5A;
		16'h4D52: out_word = 8'h46;
		16'h4D53: out_word = 8'h4A;
		16'h4D54: out_word = 8'h52;
		16'h4D55: out_word = 8'h62;
		16'h4D56: out_word = 8'h42;
		16'h4D57: out_word = 8'h00;
		16'h4D58: out_word = 8'h00;
		16'h4D59: out_word = 8'h44;
		16'h4D5A: out_word = 8'h48;
		16'h4D5B: out_word = 8'h70;
		16'h4D5C: out_word = 8'h48;
		16'h4D5D: out_word = 8'h44;
		16'h4D5E: out_word = 8'h42;
		16'h4D5F: out_word = 8'h00;
		16'h4D60: out_word = 8'h00;
		16'h4D61: out_word = 8'h1E;
		16'h4D62: out_word = 8'h22;
		16'h4D63: out_word = 8'h22;
		16'h4D64: out_word = 8'h22;
		16'h4D65: out_word = 8'h22;
		16'h4D66: out_word = 8'h42;
		16'h4D67: out_word = 8'h00;
		16'h4D68: out_word = 8'h00;
		16'h4D69: out_word = 8'h42;
		16'h4D6A: out_word = 8'h66;
		16'h4D6B: out_word = 8'h5A;
		16'h4D6C: out_word = 8'h42;
		16'h4D6D: out_word = 8'h42;
		16'h4D6E: out_word = 8'h42;
		16'h4D6F: out_word = 8'h00;
		16'h4D70: out_word = 8'h00;
		16'h4D71: out_word = 8'h42;
		16'h4D72: out_word = 8'h42;
		16'h4D73: out_word = 8'h7E;
		16'h4D74: out_word = 8'h42;
		16'h4D75: out_word = 8'h42;
		16'h4D76: out_word = 8'h42;
		16'h4D77: out_word = 8'h00;
		16'h4D78: out_word = 8'h00;
		16'h4D79: out_word = 8'h3C;
		16'h4D7A: out_word = 8'h42;
		16'h4D7B: out_word = 8'h42;
		16'h4D7C: out_word = 8'h42;
		16'h4D7D: out_word = 8'h42;
		16'h4D7E: out_word = 8'h3C;
		16'h4D7F: out_word = 8'h00;
		16'h4D80: out_word = 8'h00;
		16'h4D81: out_word = 8'h7E;
		16'h4D82: out_word = 8'h42;
		16'h4D83: out_word = 8'h42;
		16'h4D84: out_word = 8'h42;
		16'h4D85: out_word = 8'h42;
		16'h4D86: out_word = 8'h42;
		16'h4D87: out_word = 8'h00;
		16'h4D88: out_word = 8'h00;
		16'h4D89: out_word = 8'h3E;
		16'h4D8A: out_word = 8'h42;
		16'h4D8B: out_word = 8'h42;
		16'h4D8C: out_word = 8'h3E;
		16'h4D8D: out_word = 8'h22;
		16'h4D8E: out_word = 8'h42;
		16'h4D8F: out_word = 8'h00;
		16'h4D90: out_word = 8'h00;
		16'h4D91: out_word = 8'h7C;
		16'h4D92: out_word = 8'h42;
		16'h4D93: out_word = 8'h42;
		16'h4D94: out_word = 8'h7C;
		16'h4D95: out_word = 8'h40;
		16'h4D96: out_word = 8'h40;
		16'h4D97: out_word = 8'h00;
		16'h4D98: out_word = 8'h00;
		16'h4D99: out_word = 8'h3C;
		16'h4D9A: out_word = 8'h42;
		16'h4D9B: out_word = 8'h40;
		16'h4D9C: out_word = 8'h40;
		16'h4D9D: out_word = 8'h42;
		16'h4D9E: out_word = 8'h3C;
		16'h4D9F: out_word = 8'h00;
		16'h4DA0: out_word = 8'h00;
		16'h4DA1: out_word = 8'hFE;
		16'h4DA2: out_word = 8'h10;
		16'h4DA3: out_word = 8'h10;
		16'h4DA4: out_word = 8'h10;
		16'h4DA5: out_word = 8'h10;
		16'h4DA6: out_word = 8'h10;
		16'h4DA7: out_word = 8'h00;
		16'h4DA8: out_word = 8'h00;
		16'h4DA9: out_word = 8'h42;
		16'h4DAA: out_word = 8'h42;
		16'h4DAB: out_word = 8'h3E;
		16'h4DAC: out_word = 8'h02;
		16'h4DAD: out_word = 8'h42;
		16'h4DAE: out_word = 8'h3C;
		16'h4DAF: out_word = 8'h00;
		16'h4DB0: out_word = 8'h00;
		16'h4DB1: out_word = 8'h54;
		16'h4DB2: out_word = 8'h54;
		16'h4DB3: out_word = 8'h38;
		16'h4DB4: out_word = 8'h54;
		16'h4DB5: out_word = 8'h54;
		16'h4DB6: out_word = 8'h54;
		16'h4DB7: out_word = 8'h00;
		16'h4DB8: out_word = 8'h00;
		16'h4DB9: out_word = 8'h7C;
		16'h4DBA: out_word = 8'h42;
		16'h4DBB: out_word = 8'h7C;
		16'h4DBC: out_word = 8'h42;
		16'h4DBD: out_word = 8'h42;
		16'h4DBE: out_word = 8'h7C;
		16'h4DBF: out_word = 8'h00;
		16'h4DC0: out_word = 8'h00;
		16'h4DC1: out_word = 8'h40;
		16'h4DC2: out_word = 8'h40;
		16'h4DC3: out_word = 8'h7C;
		16'h4DC4: out_word = 8'h42;
		16'h4DC5: out_word = 8'h42;
		16'h4DC6: out_word = 8'h7C;
		16'h4DC7: out_word = 8'h00;
		16'h4DC8: out_word = 8'h00;
		16'h4DC9: out_word = 8'h42;
		16'h4DCA: out_word = 8'h42;
		16'h4DCB: out_word = 8'h72;
		16'h4DCC: out_word = 8'h4A;
		16'h4DCD: out_word = 8'h4A;
		16'h4DCE: out_word = 8'h72;
		16'h4DCF: out_word = 8'h00;
		16'h4DD0: out_word = 8'h00;
		16'h4DD1: out_word = 8'h3C;
		16'h4DD2: out_word = 8'h42;
		16'h4DD3: out_word = 8'h0C;
		16'h4DD4: out_word = 8'h02;
		16'h4DD5: out_word = 8'h42;
		16'h4DD6: out_word = 8'h3C;
		16'h4DD7: out_word = 8'h00;
		16'h4DD8: out_word = 8'h00;
		16'h4DD9: out_word = 8'h54;
		16'h4DDA: out_word = 8'h54;
		16'h4DDB: out_word = 8'h54;
		16'h4DDC: out_word = 8'h54;
		16'h4DDD: out_word = 8'h54;
		16'h4DDE: out_word = 8'h7C;
		16'h4DDF: out_word = 8'h00;
		16'h4DE0: out_word = 8'h00;
		16'h4DE1: out_word = 8'h3C;
		16'h4DE2: out_word = 8'h42;
		16'h4DE3: out_word = 8'h0E;
		16'h4DE4: out_word = 8'h02;
		16'h4DE5: out_word = 8'h42;
		16'h4DE6: out_word = 8'h3C;
		16'h4DE7: out_word = 8'h00;
		16'h4DE8: out_word = 8'h00;
		16'h4DE9: out_word = 8'h54;
		16'h4DEA: out_word = 8'h54;
		16'h4DEB: out_word = 8'h54;
		16'h4DEC: out_word = 8'h54;
		16'h4DED: out_word = 8'h54;
		16'h4DEE: out_word = 8'h7E;
		16'h4DEF: out_word = 8'h02;
		16'h4DF0: out_word = 8'h00;
		16'h4DF1: out_word = 8'h42;
		16'h4DF2: out_word = 8'h42;
		16'h4DF3: out_word = 8'h42;
		16'h4DF4: out_word = 8'h7E;
		16'h4DF5: out_word = 8'h02;
		16'h4DF6: out_word = 8'h02;
		16'h4DF7: out_word = 8'h00;
		16'h4DF8: out_word = 8'h3C;
		16'h4DF9: out_word = 8'h42;
		16'h4DFA: out_word = 8'h99;
		16'h4DFB: out_word = 8'hA1;
		16'h4DFC: out_word = 8'hA1;
		16'h4DFD: out_word = 8'h99;
		16'h4DFE: out_word = 8'h42;
		16'h4DFF: out_word = 8'h3C;
		16'h4E00: out_word = 8'hF3;
		16'h4E01: out_word = 8'hF5;
		16'h4E02: out_word = 8'hE5;
		16'h4E03: out_word = 8'hD5;
		16'h4E04: out_word = 8'hC5;
		16'h4E05: out_word = 8'hD9;
		16'h4E06: out_word = 8'hE5;
		16'h4E07: out_word = 8'h2A;
		16'h4E08: out_word = 8'h3D;
		16'h4E09: out_word = 8'h5C;
		16'h4E0A: out_word = 8'h22;
		16'h4E0B: out_word = 8'h32;
		16'h4E0C: out_word = 8'hF6;
		16'h4E0D: out_word = 8'h3A;
		16'h4E0E: out_word = 8'h19;
		16'h4E0F: out_word = 8'h5D;
		16'h4E10: out_word = 8'h32;
		16'h4E11: out_word = 8'hF6;
		16'h4E12: out_word = 8'h5C;
		16'h4E13: out_word = 8'hC6;
		16'h4E14: out_word = 8'h3C;
		16'h4E15: out_word = 8'h32;
		16'h4E16: out_word = 8'h16;
		16'h4E17: out_word = 8'h5D;
		16'h4E18: out_word = 8'h21;
		16'h4E19: out_word = 8'h00;
		16'h4E1A: out_word = 8'h3C;
		16'h4E1B: out_word = 8'h11;
		16'h4E1C: out_word = 8'h00;
		16'h4E1D: out_word = 8'h80;
		16'h4E1E: out_word = 8'hD5;
		16'h4E1F: out_word = 8'hED;
		16'h4E20: out_word = 8'h53;
		16'h4E21: out_word = 8'h36;
		16'h4E22: out_word = 8'h5C;
		16'h4E23: out_word = 8'h01;
		16'h4E24: out_word = 8'h00;
		16'h4E25: out_word = 8'h04;
		16'h4E26: out_word = 8'hED;
		16'h4E27: out_word = 8'hB0;
		16'h4E28: out_word = 8'hFD;
		16'h4E29: out_word = 8'h36;
		16'h4E2A: out_word = 8'h47;
		16'h4E2B: out_word = 8'h00;
		16'h4E2C: out_word = 8'hE1;
		16'h4E2D: out_word = 8'h01;
		16'h4E2E: out_word = 8'h80;
		16'h4E2F: out_word = 8'h00;
		16'h4E30: out_word = 8'hC5;
		16'h4E31: out_word = 8'h23;
		16'h4E32: out_word = 8'h23;
		16'h4E33: out_word = 8'h23;
		16'h4E34: out_word = 8'h06;
		16'h4E35: out_word = 8'h03;
		16'h4E36: out_word = 8'h56;
		16'h4E37: out_word = 8'h7A;
		16'h4E38: out_word = 8'h17;
		16'h4E39: out_word = 8'hB2;
		16'h4E3A: out_word = 8'h77;
		16'h4E3B: out_word = 8'h23;
		16'h4E3C: out_word = 8'h10;
		16'h4E3D: out_word = 8'hF8;
		16'h4E3E: out_word = 8'hC1;
		16'h4E3F: out_word = 8'h0B;
		16'h4E40: out_word = 8'h23;
		16'h4E41: out_word = 8'h23;
		16'h4E42: out_word = 8'h78;
		16'h4E43: out_word = 8'hB1;
		16'h4E44: out_word = 8'h20;
		16'h4E45: out_word = 8'hEA;
		16'h4E46: out_word = 8'hAF;
		16'h4E47: out_word = 8'hD3;
		16'h4E48: out_word = 8'hFE;
		16'h4E49: out_word = 8'h3E;
		16'h4E4A: out_word = 8'h44;
		16'h4E4B: out_word = 8'h32;
		16'h4E4C: out_word = 8'h48;
		16'h4E4D: out_word = 8'h5C;
		16'h4E4E: out_word = 8'h3D;
		16'h4E4F: out_word = 8'h3D;
		16'h4E50: out_word = 8'h32;
		16'h4E51: out_word = 8'h8D;
		16'h4E52: out_word = 8'h5C;
		16'h4E53: out_word = 8'hCD;
		16'h4E54: out_word = 8'h6B;
		16'h4E55: out_word = 8'h0D;
		16'h4E56: out_word = 8'hF3;
		16'h4E57: out_word = 8'hAF;
		16'h4E58: out_word = 8'h32;
		16'h4E59: out_word = 8'h6E;
		16'h4E5A: out_word = 8'hF8;
		16'h4E5B: out_word = 8'h21;
		16'h4E5C: out_word = 8'h09;
		16'h4E5D: out_word = 8'hFA;
		16'h4E5E: out_word = 8'hE5;
		16'h4E5F: out_word = 8'hED;
		16'h4E60: out_word = 8'h73;
		16'h4E61: out_word = 8'h3D;
		16'h4E62: out_word = 8'h5C;
		16'h4E63: out_word = 8'hFD;
		16'h4E64: out_word = 8'h36;
		16'h4E65: out_word = 8'h00;
		16'h4E66: out_word = 8'hFF;
		16'h4E67: out_word = 8'h3A;
		16'h4E68: out_word = 8'h19;
		16'h4E69: out_word = 8'h5D;
		16'h4E6A: out_word = 8'h0E;
		16'h4E6B: out_word = 8'h01;
		16'h4E6C: out_word = 8'hCD;
		16'h4E6D: out_word = 8'h13;
		16'h4E6E: out_word = 8'h3D;
		16'h4E6F: out_word = 8'h21;
		16'h4E70: out_word = 8'h00;
		16'h4E71: out_word = 8'h90;
		16'h4E72: out_word = 8'h11;
		16'h4E73: out_word = 8'h00;
		16'h4E74: out_word = 8'h00;
		16'h4E75: out_word = 8'h01;
		16'h4E76: out_word = 8'h05;
		16'h4E77: out_word = 8'h08;
		16'h4E78: out_word = 8'hCD;
		16'h4E79: out_word = 8'h13;
		16'h4E7A: out_word = 8'h3D;
		16'h4E7B: out_word = 8'hFD;
		16'h4E7C: out_word = 8'h7E;
		16'h4E7D: out_word = 8'h00;
		16'h4E7E: out_word = 8'hFE;
		16'h4E7F: out_word = 8'hFF;
		16'h4E80: out_word = 8'h20;
		16'h4E81: out_word = 8'hD4;
		16'h4E82: out_word = 8'h21;
		16'h4E83: out_word = 8'h56;
		16'h4E84: out_word = 8'hF5;
		16'h4E85: out_word = 8'h22;
		16'h4E86: out_word = 8'h5C;
		16'h4E87: out_word = 8'hF5;
		16'h4E88: out_word = 8'hD9;
		16'h4E89: out_word = 8'h11;
		16'h4E8A: out_word = 8'h00;
		16'h4E8B: out_word = 8'hA0;
		16'h4E8C: out_word = 8'hD9;
		16'h4E8D: out_word = 8'h21;
		16'h4E8E: out_word = 8'h00;
		16'h4E8F: out_word = 8'h90;
		16'h4E90: out_word = 8'h11;
		16'h4E91: out_word = 8'h08;
		16'h4E92: out_word = 8'h00;
		16'h4E93: out_word = 8'h7E;
		16'h4E94: out_word = 8'hB7;
		16'h4E95: out_word = 8'hCA;
		16'h4E96: out_word = 8'h87;
		16'h4E97: out_word = 8'hF8;
		16'h4E98: out_word = 8'h11;
		16'h4E99: out_word = 8'h08;
		16'h4E9A: out_word = 8'h00;
		16'h4E9B: out_word = 8'h19;
		16'h4E9C: out_word = 8'h7E;
		16'h4E9D: out_word = 8'hFE;
		16'h4E9E: out_word = 8'h42;
		16'h4E9F: out_word = 8'hCC;
		16'h4EA0: out_word = 8'h36;
		16'h4EA1: out_word = 8'hF8;
		16'h4EA2: out_word = 8'h19;
		16'h4EA3: out_word = 8'h7E;
		16'h4EA4: out_word = 8'hB7;
		16'h4EA5: out_word = 8'h20;
		16'h4EA6: out_word = 8'hF1;
		16'h4EA7: out_word = 8'h3A;
		16'h4EA8: out_word = 8'h6E;
		16'h4EA9: out_word = 8'hF8;
		16'h4EAA: out_word = 8'hB7;
		16'h4EAB: out_word = 8'hCA;
		16'h4EAC: out_word = 8'h87;
		16'h4EAD: out_word = 8'hF8;
		16'h4EAE: out_word = 8'h06;
		16'h4EAF: out_word = 8'h3F;
		16'h4EB0: out_word = 8'h98;
		16'h4EB1: out_word = 8'hD2;
		16'h4EB2: out_word = 8'hA6;
		16'h4EB3: out_word = 8'hF8;
		16'h4EB4: out_word = 8'h3A;
		16'h4EB5: out_word = 8'h6E;
		16'h4EB6: out_word = 8'hF8;
		16'h4EB7: out_word = 8'h3D;
		16'h4EB8: out_word = 8'h32;
		16'h4EB9: out_word = 8'h6F;
		16'h4EBA: out_word = 8'hF8;
		16'h4EBB: out_word = 8'hCD;
		16'h4EBC: out_word = 8'hBB;
		16'h4EBD: out_word = 8'hF9;
		16'h4EBE: out_word = 8'h32;
		16'h4EBF: out_word = 8'h53;
		16'h4EC0: out_word = 8'hF6;
		16'h4EC1: out_word = 8'hCD;
		16'h4EC2: out_word = 8'h6B;
		16'h4EC3: out_word = 8'h0D;
		16'h4EC4: out_word = 8'hF3;
		16'h4EC5: out_word = 8'hCD;
		16'h4EC6: out_word = 8'h70;
		16'h4EC7: out_word = 8'hF8;
		16'h4EC8: out_word = 8'h3E;
		16'h4EC9: out_word = 8'h02;
		16'h4ECA: out_word = 8'hCD;
		16'h4ECB: out_word = 8'hCB;
		16'h4ECC: out_word = 8'hF8;
		16'h4ECD: out_word = 8'h3E;
		16'h4ECE: out_word = 8'h02;
		16'h4ECF: out_word = 8'hCD;
		16'h4ED0: out_word = 8'h01;
		16'h4ED1: out_word = 8'h16;
		16'h4ED2: out_word = 8'hFD;
		16'h4ED3: out_word = 8'h36;
		16'h4ED4: out_word = 8'h47;
		16'h4ED5: out_word = 8'h00;
		16'h4ED6: out_word = 8'h11;
		16'h4ED7: out_word = 8'h00;
		16'h4ED8: out_word = 8'hA0;
		16'h4ED9: out_word = 8'h21;
		16'h4EDA: out_word = 8'h08;
		16'h4EDB: out_word = 8'h00;
		16'h4EDC: out_word = 8'h3E;
		16'h4EDD: out_word = 8'h20;
		16'h4EDE: out_word = 8'hD7;
		16'h4EDF: out_word = 8'h3E;
		16'h4EE0: out_word = 8'h20;
		16'h4EE1: out_word = 8'hD7;
		16'h4EE2: out_word = 8'h01;
		16'h4EE3: out_word = 8'h08;
		16'h4EE4: out_word = 8'h00;
		16'h4EE5: out_word = 8'hD5;
		16'h4EE6: out_word = 8'hCD;
		16'h4EE7: out_word = 8'h3C;
		16'h4EE8: out_word = 8'h20;
		16'h4EE9: out_word = 8'hD1;
		16'h4EEA: out_word = 8'hEB;
		16'h4EEB: out_word = 8'hED;
		16'h4EEC: out_word = 8'h5A;
		16'h4EED: out_word = 8'hEB;
		16'h4EEE: out_word = 8'h3A;
		16'h4EEF: out_word = 8'h6E;
		16'h4EF0: out_word = 8'hF8;
		16'h4EF1: out_word = 8'h3D;
		16'h4EF2: out_word = 8'h32;
		16'h4EF3: out_word = 8'h6E;
		16'h4EF4: out_word = 8'hF8;
		16'h4EF5: out_word = 8'h28;
		16'h4EF6: out_word = 8'h3E;
		16'h4EF7: out_word = 8'h3E;
		16'h4EF8: out_word = 8'h20;
		16'h4EF9: out_word = 8'hD7;
		16'h4EFA: out_word = 8'h3E;
		16'h4EFB: out_word = 8'h20;
		16'h4EFC: out_word = 8'hD7;
		16'h4EFD: out_word = 8'h01;
		16'h4EFE: out_word = 8'h08;
		16'h4EFF: out_word = 8'h00;
		16'h4F00: out_word = 8'hD5;
		16'h4F01: out_word = 8'hCD;
		16'h4F02: out_word = 8'h3C;
		16'h4F03: out_word = 8'h20;
		16'h4F04: out_word = 8'hD1;
		16'h4F05: out_word = 8'hEB;
		16'h4F06: out_word = 8'hED;
		16'h4F07: out_word = 8'h5A;
		16'h4F08: out_word = 8'hEB;
		16'h4F09: out_word = 8'h3A;
		16'h4F0A: out_word = 8'h6E;
		16'h4F0B: out_word = 8'hF8;
		16'h4F0C: out_word = 8'h3D;
		16'h4F0D: out_word = 8'h32;
		16'h4F0E: out_word = 8'h6E;
		16'h4F0F: out_word = 8'hF8;
		16'h4F10: out_word = 8'h28;
		16'h4F11: out_word = 8'h23;
		16'h4F12: out_word = 8'h3E;
		16'h4F13: out_word = 8'h20;
		16'h4F14: out_word = 8'hD7;
		16'h4F15: out_word = 8'h3E;
		16'h4F16: out_word = 8'h20;
		16'h4F17: out_word = 8'hD7;
		16'h4F18: out_word = 8'h01;
		16'h4F19: out_word = 8'h08;
		16'h4F1A: out_word = 8'h00;
		16'h4F1B: out_word = 8'hD5;
		16'h4F1C: out_word = 8'hCD;
		16'h4F1D: out_word = 8'h3C;
		16'h4F1E: out_word = 8'h20;
		16'h4F1F: out_word = 8'hD1;
		16'h4F20: out_word = 8'hEB;
		16'h4F21: out_word = 8'hED;
		16'h4F22: out_word = 8'h5A;
		16'h4F23: out_word = 8'hEB;
		16'h4F24: out_word = 8'h3A;
		16'h4F25: out_word = 8'h6E;
		16'h4F26: out_word = 8'hF8;
		16'h4F27: out_word = 8'h3D;
		16'h4F28: out_word = 8'h32;
		16'h4F29: out_word = 8'h6E;
		16'h4F2A: out_word = 8'hF8;
		16'h4F2B: out_word = 8'h28;
		16'h4F2C: out_word = 8'h08;
		16'h4F2D: out_word = 8'h3E;
		16'h4F2E: out_word = 8'h06;
		16'h4F2F: out_word = 8'hD7;
		16'h4F30: out_word = 8'h18;
		16'h4F31: out_word = 8'hAA;
		16'h4F32: out_word = 8'h00;
		16'h4F33: out_word = 8'h00;
		16'h4F34: out_word = 8'h00;
		16'h4F35: out_word = 8'h21;
		16'h4F36: out_word = 8'h02;
		16'h4F37: out_word = 8'h58;
		16'h4F38: out_word = 8'hCD;
		16'h4F39: out_word = 8'h16;
		16'h4F3A: out_word = 8'hF8;
		16'h4F3B: out_word = 8'h11;
		16'h4F3C: out_word = 8'h0A;
		16'h4F3D: out_word = 8'h00;
		16'h4F3E: out_word = 8'hDD;
		16'h4F3F: out_word = 8'h21;
		16'h4F40: out_word = 8'h34;
		16'h4F41: out_word = 8'hF6;
		16'h4F42: out_word = 8'hDD;
		16'h4F43: out_word = 8'h36;
		16'h4F44: out_word = 8'h00;
		16'h4F45: out_word = 8'h00;
		16'h4F46: out_word = 8'hFB;
		16'h4F47: out_word = 8'hFD;
		16'h4F48: out_word = 8'hCB;
		16'h4F49: out_word = 8'h01;
		16'h4F4A: out_word = 8'hAE;
		16'h4F4B: out_word = 8'h76;
		16'h4F4C: out_word = 8'hE5;
		16'h4F4D: out_word = 8'hDD;
		16'h4F4E: out_word = 8'hE5;
		16'h4F4F: out_word = 8'hCD;
		16'h4F50: out_word = 8'hBB;
		16'h4F51: out_word = 8'hF9;
		16'h4F52: out_word = 8'hFE;
		16'h4F53: out_word = 8'h40;
		16'h4F54: out_word = 8'hC2;
		16'h4F55: out_word = 8'h92;
		16'h4F56: out_word = 8'hF7;
		16'h4F57: out_word = 8'hCD;
		16'h4F58: out_word = 8'h89;
		16'h4F59: out_word = 8'hF9;
		16'h4F5A: out_word = 8'hDD;
		16'h4F5B: out_word = 8'hE1;
		16'h4F5C: out_word = 8'hE1;
		16'h4F5D: out_word = 8'hFD;
		16'h4F5E: out_word = 8'hCB;
		16'h4F5F: out_word = 8'h01;
		16'h4F60: out_word = 8'h6E;
		16'h4F61: out_word = 8'h28;
		16'h4F62: out_word = 8'hE3;
		16'h4F63: out_word = 8'h3A;
		16'h4F64: out_word = 8'h08;
		16'h4F65: out_word = 8'h5C;
		16'h4F66: out_word = 8'hFE;
		16'h4F67: out_word = 8'h08;
		16'h4F68: out_word = 8'hCA;
		16'h4F69: out_word = 8'hED;
		16'h4F6A: out_word = 8'hF6;
		16'h4F6B: out_word = 8'hFE;
		16'h4F6C: out_word = 8'h6F;
		16'h4F6D: out_word = 8'h28;
		16'h4F6E: out_word = 8'h7E;
		16'h4F6F: out_word = 8'hFE;
		16'h4F70: out_word = 8'h36;
		16'h4F71: out_word = 8'h28;
		16'h4F72: out_word = 8'h7A;
		16'h4F73: out_word = 8'hFE;
		16'h4F74: out_word = 8'h09;
		16'h4F75: out_word = 8'hCA;
		16'h4F76: out_word = 8'h0C;
		16'h4F77: out_word = 8'hF7;
		16'h4F78: out_word = 8'hFE;
		16'h4F79: out_word = 8'h70;
		16'h4F7A: out_word = 8'hCA;
		16'h4F7B: out_word = 8'h0C;
		16'h4F7C: out_word = 8'hF7;
		16'h4F7D: out_word = 8'hFE;
		16'h4F7E: out_word = 8'h37;
		16'h4F7F: out_word = 8'hCA;
		16'h4F80: out_word = 8'h0C;
		16'h4F81: out_word = 8'hF7;
		16'h4F82: out_word = 8'hFE;
		16'h4F83: out_word = 8'h0B;
		16'h4F84: out_word = 8'hCA;
		16'h4F85: out_word = 8'h2E;
		16'h4F86: out_word = 8'hF7;
		16'h4F87: out_word = 8'hFE;
		16'h4F88: out_word = 8'h71;
		16'h4F89: out_word = 8'hCA;
		16'h4F8A: out_word = 8'h2E;
		16'h4F8B: out_word = 8'hF7;
		16'h4F8C: out_word = 8'hFE;
		16'h4F8D: out_word = 8'h39;
		16'h4F8E: out_word = 8'hCA;
		16'h4F8F: out_word = 8'h2E;
		16'h4F90: out_word = 8'hF7;
		16'h4F91: out_word = 8'hFE;
		16'h4F92: out_word = 8'h0A;
		16'h4F93: out_word = 8'hCA;
		16'h4F94: out_word = 8'h64;
		16'h4F95: out_word = 8'hF7;
		16'h4F96: out_word = 8'hFE;
		16'h4F97: out_word = 8'h61;
		16'h4F98: out_word = 8'hCA;
		16'h4F99: out_word = 8'h64;
		16'h4F9A: out_word = 8'hF7;
		16'h4F9B: out_word = 8'hFE;
		16'h4F9C: out_word = 8'h38;
		16'h4F9D: out_word = 8'hCA;
		16'h4F9E: out_word = 8'h64;
		16'h4F9F: out_word = 8'hF7;
		16'h4FA0: out_word = 8'hFE;
		16'h4FA1: out_word = 8'h64;
		16'h4FA2: out_word = 8'hCA;
		16'h4FA3: out_word = 8'h1B;
		16'h4FA4: out_word = 8'hFA;
		16'h4FA5: out_word = 8'hFE;
		16'h4FA6: out_word = 8'h31;
		16'h4FA7: out_word = 8'h28;
		16'h4FA8: out_word = 8'h27;
		16'h4FA9: out_word = 8'hFE;
		16'h4FAA: out_word = 8'h32;
		16'h4FAB: out_word = 8'h28;
		16'h4FAC: out_word = 8'h23;
		16'h4FAD: out_word = 8'hFE;
		16'h4FAE: out_word = 8'h33;
		16'h4FAF: out_word = 8'h28;
		16'h4FB0: out_word = 8'h1F;
		16'h4FB1: out_word = 8'hFE;
		16'h4FB2: out_word = 8'h34;
		16'h4FB3: out_word = 8'h28;
		16'h4FB4: out_word = 8'h1B;
		16'h4FB5: out_word = 8'hF5;
		16'h4FB6: out_word = 8'h3E;
		16'h4FB7: out_word = 8'hFE;
		16'h4FB8: out_word = 8'hDB;
		16'h4FB9: out_word = 8'hFE;
		16'h4FBA: out_word = 8'h1F;
		16'h4FBB: out_word = 8'h30;
		16'h4FBC: out_word = 8'h89;
		16'h4FBD: out_word = 8'hF1;
		16'h4FBE: out_word = 8'hFE;
		16'h4FBF: out_word = 8'h0D;
		16'h4FC0: out_word = 8'hCA;
		16'h4FC1: out_word = 8'h9D;
		16'h4FC2: out_word = 8'hF7;
		16'h4FC3: out_word = 8'hFE;
		16'h4FC4: out_word = 8'h30;
		16'h4FC5: out_word = 8'hCA;
		16'h4FC6: out_word = 8'h9D;
		16'h4FC7: out_word = 8'hF7;
		16'h4FC8: out_word = 8'hFE;
		16'h4FC9: out_word = 8'h20;
		16'h4FCA: out_word = 8'hCA;
		16'h4FCB: out_word = 8'h9D;
		16'h4FCC: out_word = 8'hF7;
		16'h4FCD: out_word = 8'hC3;
		16'h4FCE: out_word = 8'h46;
		16'h4FCF: out_word = 8'hF6;
		16'h4FD0: out_word = 8'hF5;
		16'h4FD1: out_word = 8'hCD;
		16'h4FD2: out_word = 8'h6B;
		16'h4FD3: out_word = 8'h0D;
		16'h4FD4: out_word = 8'h3E;
		16'h4FD5: out_word = 8'h03;
		16'h4FD6: out_word = 8'hCD;
		16'h4FD7: out_word = 8'hCB;
		16'h4FD8: out_word = 8'hF8;
		16'h4FD9: out_word = 8'hF1;
		16'h4FDA: out_word = 8'hD6;
		16'h4FDB: out_word = 8'h31;
		16'h4FDC: out_word = 8'h0E;
		16'h4FDD: out_word = 8'h01;
		16'h4FDE: out_word = 8'h32;
		16'h4FDF: out_word = 8'hF8;
		16'h4FE0: out_word = 8'h5C;
		16'h4FE1: out_word = 8'h32;
		16'h4FE2: out_word = 8'hF9;
		16'h4FE3: out_word = 8'h5C;
		16'h4FE4: out_word = 8'h32;
		16'h4FE5: out_word = 8'h19;
		16'h4FE6: out_word = 8'h5D;
		16'h4FE7: out_word = 8'hCD;
		16'h4FE8: out_word = 8'h13;
		16'h4FE9: out_word = 8'h3D;
		16'h4FEA: out_word = 8'hC3;
		16'h4FEB: out_word = 8'h56;
		16'h4FEC: out_word = 8'hF5;
		16'h4FED: out_word = 8'hCD;
		16'h4FEE: out_word = 8'h70;
		16'h4FEF: out_word = 8'hF8;
		16'h4FF0: out_word = 8'hCD;
		16'h4FF1: out_word = 8'h26;
		16'h4FF2: out_word = 8'hF8;
		16'h4FF3: out_word = 8'hDD;
		16'h4FF4: out_word = 8'h35;
		16'h4FF5: out_word = 8'hFF;
		16'h4FF6: out_word = 8'hFF;
		16'h4FF7: out_word = 8'hFF;
		16'h4FF8: out_word = 8'hFF;
		16'h4FF9: out_word = 8'hFF;
		16'h4FFA: out_word = 8'hFF;
		16'h4FFB: out_word = 8'hFF;
		16'h4FFC: out_word = 8'hFF;
		16'h4FFD: out_word = 8'hFF;
		16'h4FFE: out_word = 8'hFF;
		16'h4FFF: out_word = 8'hFF;
		16'h5000: out_word = 8'h16;
		16'h5001: out_word = 8'h09;
		16'h5002: out_word = 8'h05;
		16'h5003: out_word = 8'h46;
		16'h5004: out_word = 8'h6F;
		16'h5005: out_word = 8'h75;
		16'h5006: out_word = 8'h6E;
		16'h5007: out_word = 8'h64;
		16'h5008: out_word = 8'h20;
		16'h5009: out_word = 8'h52;
		16'h500A: out_word = 8'h41;
		16'h500B: out_word = 8'h4D;
		16'h500C: out_word = 8'h44;
		16'h500D: out_word = 8'h49;
		16'h500E: out_word = 8'h53;
		16'h500F: out_word = 8'h4B;
		16'h5010: out_word = 8'h20;
		16'h5011: out_word = 8'h6D;
		16'h5012: out_word = 8'h65;
		16'h5013: out_word = 8'h6D;
		16'h5014: out_word = 8'h6F;
		16'h5015: out_word = 8'h72;
		16'h5016: out_word = 8'h79;
		16'h5017: out_word = 8'h00;
		16'h5018: out_word = 8'hCD;
		16'h5019: out_word = 8'hDF;
		16'h501A: out_word = 8'h1D;
		16'h501B: out_word = 8'hCD;
		16'h501C: out_word = 8'h75;
		16'h501D: out_word = 8'h1D;
		16'h501E: out_word = 8'hCD;
		16'h501F: out_word = 8'h31;
		16'h5020: out_word = 8'h05;
		16'h5021: out_word = 8'h1A;
		16'h5022: out_word = 8'hCD;
		16'h5023: out_word = 8'h24;
		16'h5024: out_word = 8'h05;
		16'h5025: out_word = 8'h32;
		16'h5026: out_word = 8'h19;
		16'h5027: out_word = 8'h5D;
		16'h5028: out_word = 8'hCD;
		16'h5029: out_word = 8'hCB;
		16'h502A: out_word = 8'h3D;
		16'h502B: out_word = 8'hC3;
		16'h502C: out_word = 8'hE1;
		16'h502D: out_word = 8'h03;
		16'h502E: out_word = 8'h06;
		16'h502F: out_word = 8'h43;
		16'h5030: out_word = 8'h3A;
		16'h5031: out_word = 8'hD6;
		16'h5032: out_word = 8'h5C;
		16'h5033: out_word = 8'hB7;
		16'h5034: out_word = 8'h20;
		16'h5035: out_word = 8'h17;
		16'h5036: out_word = 8'hCD;
		16'h5037: out_word = 8'h8C;
		16'h5038: out_word = 8'h1D;
		16'h5039: out_word = 8'hFE;
		16'h503A: out_word = 8'hAF;
		16'h503B: out_word = 8'h06;
		16'h503C: out_word = 8'h43;
		16'h503D: out_word = 8'h28;
		16'h503E: out_word = 8'h0E;
		16'h503F: out_word = 8'hFE;
		16'h5040: out_word = 8'hE4;
		16'h5041: out_word = 8'h06;
		16'h5042: out_word = 8'h44;
		16'h5043: out_word = 8'h28;
		16'h5044: out_word = 8'h08;
		16'h5045: out_word = 8'hFE;
		16'h5046: out_word = 8'h23;
		16'h5047: out_word = 8'h06;
		16'h5048: out_word = 8'h23;
		16'h5049: out_word = 8'h28;
		16'h504A: out_word = 8'h02;
		16'h504B: out_word = 8'h06;
		16'h504C: out_word = 8'h42;
		16'h504D: out_word = 8'h21;
		16'h504E: out_word = 8'hE5;
		16'h504F: out_word = 8'h5C;
		16'h5050: out_word = 8'h70;
		16'h5051: out_word = 8'hC9;
		16'h5052: out_word = 8'hF3;
		16'h5053: out_word = 8'hE5;
		16'h5054: out_word = 8'hC5;
		16'h5055: out_word = 8'hD5;
		16'h5056: out_word = 8'hE7;
		16'h5057: out_word = 8'h8E;
		16'h5058: out_word = 8'h02;
		16'h5059: out_word = 8'h0E;
		16'h505A: out_word = 8'h00;
		16'h505B: out_word = 8'h20;
		16'h505C: out_word = 8'hF9;
		16'h505D: out_word = 8'hE7;
		16'h505E: out_word = 8'h1E;
		16'h505F: out_word = 8'h03;
		16'h5060: out_word = 8'h30;
		16'h5061: out_word = 8'hF4;
		16'h5062: out_word = 8'h15;
		16'h5063: out_word = 8'h5F;
		16'h5064: out_word = 8'hE7;
		16'h5065: out_word = 8'h33;
		16'h5066: out_word = 8'h03;
		16'h5067: out_word = 8'hD1;
		16'h5068: out_word = 8'hC1;
		16'h5069: out_word = 8'hE1;
		16'h506A: out_word = 8'hE6;
		16'h506B: out_word = 8'hDF;
		16'h506C: out_word = 8'hFB;
		16'h506D: out_word = 8'hC9;
		16'h506E: out_word = 8'h21;
		16'h506F: out_word = 8'hE5;
		16'h5070: out_word = 8'h58;
		16'h5071: out_word = 8'h06;
		16'h5072: out_word = 8'h0A;
		16'h5073: out_word = 8'h36;
		16'h5074: out_word = 8'h07;
		16'h5075: out_word = 8'h23;
		16'h5076: out_word = 8'h10;
		16'h5077: out_word = 8'hFB;
		16'h5078: out_word = 8'h36;
		16'h5079: out_word = 8'h02;
		16'h507A: out_word = 8'h23;
		16'h507B: out_word = 8'h36;
		16'h507C: out_word = 8'h16;
		16'h507D: out_word = 8'h23;
		16'h507E: out_word = 8'h36;
		16'h507F: out_word = 8'h34;
		16'h5080: out_word = 8'h23;
		16'h5081: out_word = 8'h36;
		16'h5082: out_word = 8'h25;
		16'h5083: out_word = 8'h23;
		16'h5084: out_word = 8'h36;
		16'h5085: out_word = 8'h28;
		16'h5086: out_word = 8'h23;
		16'h5087: out_word = 8'h36;
		16'h5088: out_word = 8'h07;
		16'h5089: out_word = 8'h21;
		16'h508A: out_word = 8'hEE;
		16'h508B: out_word = 8'h40;
		16'h508C: out_word = 8'h06;
		16'h508D: out_word = 8'h08;
		16'h508E: out_word = 8'hAF;
		16'h508F: out_word = 8'hC5;
		16'h5090: out_word = 8'h37;
		16'h5091: out_word = 8'h17;
		16'h5092: out_word = 8'hE5;
		16'h5093: out_word = 8'hF5;
		16'h5094: out_word = 8'h06;
		16'h5095: out_word = 8'h05;
		16'h5096: out_word = 8'h23;
		16'h5097: out_word = 8'h77;
		16'h5098: out_word = 8'h10;
		16'h5099: out_word = 8'hFC;
		16'h509A: out_word = 8'hF1;
		16'h509B: out_word = 8'hE1;
		16'h509C: out_word = 8'hC1;
		16'h509D: out_word = 8'h11;
		16'h509E: out_word = 8'h00;
		16'h509F: out_word = 8'h01;
		16'h50A0: out_word = 8'h19;
		16'h50A1: out_word = 8'h10;
		16'h50A2: out_word = 8'hEC;
		16'h50A3: out_word = 8'hC9;
		16'h50A4: out_word = 8'hC9;
		16'h50A5: out_word = 8'h20;
		16'h50A6: out_word = 8'h44;
		16'h50A7: out_word = 8'h65;
		16'h50A8: out_word = 8'h6C;
		16'h50A9: out_word = 8'h2E;
		16'h50AA: out_word = 8'h20;
		16'h50AB: out_word = 8'h46;
		16'h50AC: out_word = 8'h69;
		16'h50AD: out_word = 8'h6C;
		16'h50AE: out_word = 8'h65;
		16'h50AF: out_word = 8'h28;
		16'h50B0: out_word = 8'h73;
		16'h50B1: out_word = 8'h29;
		16'h50B2: out_word = 8'h00;
		16'h50B3: out_word = 8'h54;
		16'h50B4: out_word = 8'h69;
		16'h50B5: out_word = 8'h74;
		16'h50B6: out_word = 8'h6C;
		16'h50B7: out_word = 8'h65;
		16'h50B8: out_word = 8'h3A;
		16'h50B9: out_word = 8'hA0;
		16'h50BA: out_word = 8'h17;
		16'h50BB: out_word = 8'h11;
		16'h50BC: out_word = 8'h20;
		16'h50BD: out_word = 8'h44;
		16'h50BE: out_word = 8'h69;
		16'h50BF: out_word = 8'h73;
		16'h50C0: out_word = 8'h6B;
		16'h50C1: out_word = 8'h20;
		16'h50C2: out_word = 8'h44;
		16'h50C3: out_word = 8'h72;
		16'h50C4: out_word = 8'h69;
		16'h50C5: out_word = 8'h76;
		16'h50C6: out_word = 8'h65;
		16'h50C7: out_word = 8'h3A;
		16'h50C8: out_word = 8'h20;
		16'h50C9: out_word = 8'h00;
		16'h50CA: out_word = 8'h17;
		16'h50CB: out_word = 8'h10;
		16'h50CC: out_word = 8'h20;
		16'h50CD: out_word = 8'h00;
		16'h50CE: out_word = 8'h17;
		16'h50CF: out_word = 8'h10;
		16'h50D0: out_word = 8'h20;
		16'h50D1: out_word = 8'h34;
		16'h50D2: out_word = 8'h30;
		16'h50D3: out_word = 8'h20;
		16'h50D4: out_word = 8'h54;
		16'h50D5: out_word = 8'h72;
		16'h50D6: out_word = 8'h61;
		16'h50D7: out_word = 8'h63;
		16'h50D8: out_word = 8'h6B;
		16'h50D9: out_word = 8'h20;
		16'h50DA: out_word = 8'h53;
		16'h50DB: out_word = 8'h2E;
		16'h50DC: out_word = 8'h20;
		16'h50DD: out_word = 8'h53;
		16'h50DE: out_word = 8'h69;
		16'h50DF: out_word = 8'h64;
		16'h50E0: out_word = 8'h65;
		16'h50E1: out_word = 8'h00;
		16'h50E2: out_word = 8'h17;
		16'h50E3: out_word = 8'h10;
		16'h50E4: out_word = 8'h20;
		16'h50E5: out_word = 8'h38;
		16'h50E6: out_word = 8'h30;
		16'h50E7: out_word = 8'h20;
		16'h50E8: out_word = 8'h54;
		16'h50E9: out_word = 8'h72;
		16'h50EA: out_word = 8'h61;
		16'h50EB: out_word = 8'h63;
		16'h50EC: out_word = 8'h6B;
		16'h50ED: out_word = 8'h20;
		16'h50EE: out_word = 8'h53;
		16'h50EF: out_word = 8'h2E;
		16'h50F0: out_word = 8'h20;
		16'h50F1: out_word = 8'h53;
		16'h50F2: out_word = 8'h69;
		16'h50F3: out_word = 8'h64;
		16'h50F4: out_word = 8'h65;
		16'h50F5: out_word = 8'h00;
		16'h50F6: out_word = 8'h17;
		16'h50F7: out_word = 8'h10;
		16'h50F8: out_word = 8'h20;
		16'h50F9: out_word = 8'h34;
		16'h50FA: out_word = 8'h30;
		16'h50FB: out_word = 8'h20;
		16'h50FC: out_word = 8'h54;
		16'h50FD: out_word = 8'h72;
		16'h50FE: out_word = 8'h61;
		16'h50FF: out_word = 8'h63;
		16'h5100: out_word = 8'h6B;
		16'h5101: out_word = 8'h20;
		16'h5102: out_word = 8'h44;
		16'h5103: out_word = 8'h2E;
		16'h5104: out_word = 8'h20;
		16'h5105: out_word = 8'h53;
		16'h5106: out_word = 8'h69;
		16'h5107: out_word = 8'h64;
		16'h5108: out_word = 8'h65;
		16'h5109: out_word = 8'h00;
		16'h510A: out_word = 8'h17;
		16'h510B: out_word = 8'h10;
		16'h510C: out_word = 8'h20;
		16'h510D: out_word = 8'h38;
		16'h510E: out_word = 8'h30;
		16'h510F: out_word = 8'h20;
		16'h5110: out_word = 8'h54;
		16'h5111: out_word = 8'h72;
		16'h5112: out_word = 8'h61;
		16'h5113: out_word = 8'h63;
		16'h5114: out_word = 8'h6B;
		16'h5115: out_word = 8'h20;
		16'h5116: out_word = 8'h44;
		16'h5117: out_word = 8'h2E;
		16'h5118: out_word = 8'h20;
		16'h5119: out_word = 8'h53;
		16'h511A: out_word = 8'h69;
		16'h511B: out_word = 8'h64;
		16'h511C: out_word = 8'h65;
		16'h511D: out_word = 8'h00;
		16'h511E: out_word = 8'h17;
		16'h511F: out_word = 8'h10;
		16'h5120: out_word = 8'h20;
		16'h5121: out_word = 8'h46;
		16'h5122: out_word = 8'h72;
		16'h5123: out_word = 8'h65;
		16'h5124: out_word = 8'h65;
		16'h5125: out_word = 8'h20;
		16'h5126: out_word = 8'h53;
		16'h5127: out_word = 8'h65;
		16'h5128: out_word = 8'h63;
		16'h5129: out_word = 8'h74;
		16'h512A: out_word = 8'h6F;
		16'h512B: out_word = 8'h72;
		16'h512C: out_word = 8'h20;
		16'h512D: out_word = 8'h00;
		16'h512E: out_word = 8'h0D;
		16'h512F: out_word = 8'h0D;
		16'h5130: out_word = 8'h20;
		16'h5131: out_word = 8'h20;
		16'h5132: out_word = 8'h46;
		16'h5133: out_word = 8'h69;
		16'h5134: out_word = 8'h6C;
		16'h5135: out_word = 8'h65;
		16'h5136: out_word = 8'h20;
		16'h5137: out_word = 8'h4E;
		16'h5138: out_word = 8'h61;
		16'h5139: out_word = 8'h6D;
		16'h513A: out_word = 8'h65;
		16'h513B: out_word = 8'h20;
		16'h513C: out_word = 8'h20;
		16'h513D: out_word = 8'h20;
		16'h513E: out_word = 8'h20;
		16'h513F: out_word = 8'h53;
		16'h5140: out_word = 8'h74;
		16'h5141: out_word = 8'h61;
		16'h5142: out_word = 8'h72;
		16'h5143: out_word = 8'h74;
		16'h5144: out_word = 8'h20;
		16'h5145: out_word = 8'h4C;
		16'h5146: out_word = 8'h65;
		16'h5147: out_word = 8'h6E;
		16'h5148: out_word = 8'h67;
		16'h5149: out_word = 8'h74;
		16'h514A: out_word = 8'h68;
		16'h514B: out_word = 8'h20;
		16'h514C: out_word = 8'h4C;
		16'h514D: out_word = 8'h69;
		16'h514E: out_word = 8'h6E;
		16'h514F: out_word = 8'h65;
		16'h5150: out_word = 8'h00;
		16'h5151: out_word = 8'h2A;
		16'h5152: out_word = 8'h61;
		16'h5153: out_word = 8'h5C;
		16'h5154: out_word = 8'h22;
		16'h5155: out_word = 8'hCF;
		16'h5156: out_word = 8'h5C;
		16'h5157: out_word = 8'h01;
		16'h5158: out_word = 8'h22;
		16'h5159: out_word = 8'h02;
		16'h515A: out_word = 8'hC3;
		16'h515B: out_word = 8'h23;
		16'h515C: out_word = 8'h1E;
		16'h515D: out_word = 8'hAF;
		16'h515E: out_word = 8'h11;
		16'h515F: out_word = 8'h10;
		16'h5160: out_word = 8'h27;
		16'h5161: out_word = 8'hED;
		16'h5162: out_word = 8'h52;
		16'h5163: out_word = 8'h38;
		16'h5164: out_word = 8'h03;
		16'h5165: out_word = 8'h3C;
		16'h5166: out_word = 8'h18;
		16'h5167: out_word = 8'hF9;
		16'h5168: out_word = 8'hC6;
		16'h5169: out_word = 8'h30;
		16'h516A: out_word = 8'hCD;
		16'h516B: out_word = 8'hA8;
		16'h516C: out_word = 8'h11;
		16'h516D: out_word = 8'h19;
		16'h516E: out_word = 8'hAF;
		16'h516F: out_word = 8'h11;
		16'h5170: out_word = 8'hE8;
		16'h5171: out_word = 8'h03;
		16'h5172: out_word = 8'hED;
		16'h5173: out_word = 8'h52;
		16'h5174: out_word = 8'h38;
		16'h5175: out_word = 8'h03;
		16'h5176: out_word = 8'h3C;
		16'h5177: out_word = 8'h18;
		16'h5178: out_word = 8'hF9;
		16'h5179: out_word = 8'hC6;
		16'h517A: out_word = 8'h30;
		16'h517B: out_word = 8'hCD;
		16'h517C: out_word = 8'hA8;
		16'h517D: out_word = 8'h11;
		16'h517E: out_word = 8'h19;
		16'h517F: out_word = 8'hAF;
		16'h5180: out_word = 8'h11;
		16'h5181: out_word = 8'h64;
		16'h5182: out_word = 8'h00;
		16'h5183: out_word = 8'hED;
		16'h5184: out_word = 8'h52;
		16'h5185: out_word = 8'h38;
		16'h5186: out_word = 8'h03;
		16'h5187: out_word = 8'h3C;
		16'h5188: out_word = 8'h18;
		16'h5189: out_word = 8'hF9;
		16'h518A: out_word = 8'hC6;
		16'h518B: out_word = 8'h30;
		16'h518C: out_word = 8'hCD;
		16'h518D: out_word = 8'hA8;
		16'h518E: out_word = 8'h11;
		16'h518F: out_word = 8'h19;
		16'h5190: out_word = 8'hAF;
		16'h5191: out_word = 8'h11;
		16'h5192: out_word = 8'h0A;
		16'h5193: out_word = 8'h00;
		16'h5194: out_word = 8'hED;
		16'h5195: out_word = 8'h52;
		16'h5196: out_word = 8'h38;
		16'h5197: out_word = 8'h03;
		16'h5198: out_word = 8'h3C;
		16'h5199: out_word = 8'h18;
		16'h519A: out_word = 8'hF9;
		16'h519B: out_word = 8'hC6;
		16'h519C: out_word = 8'h30;
		16'h519D: out_word = 8'hCD;
		16'h519E: out_word = 8'hA8;
		16'h519F: out_word = 8'h11;
		16'h51A0: out_word = 8'h19;
		16'h51A1: out_word = 8'h7D;
		16'h51A2: out_word = 8'hC6;
		16'h51A3: out_word = 8'h30;
		16'h51A4: out_word = 8'hCD;
		16'h51A5: out_word = 8'hA8;
		16'h51A6: out_word = 8'h11;
		16'h51A7: out_word = 8'hC9;
		16'h51A8: out_word = 8'hE5;
		16'h51A9: out_word = 8'hD5;
		16'h51AA: out_word = 8'hCD;
		16'h51AB: out_word = 8'h82;
		16'h51AC: out_word = 8'h3D;
		16'h51AD: out_word = 8'hD1;
		16'h51AE: out_word = 8'hE1;
		16'h51AF: out_word = 8'hC9;
		16'h51B0: out_word = 8'hE5;
		16'h51B1: out_word = 8'hC5;
		16'h51B2: out_word = 8'h3A;
		16'h51B3: out_word = 8'hF9;
		16'h51B4: out_word = 8'h5C;
		16'h51B5: out_word = 8'h21;
		16'h51B6: out_word = 8'hF6;
		16'h51B7: out_word = 8'h5C;
		16'h51B8: out_word = 8'hBE;
		16'h51B9: out_word = 8'hC4;
		16'h51BA: out_word = 8'hCB;
		16'h51BB: out_word = 8'h3D;
		16'h51BC: out_word = 8'hC1;
		16'h51BD: out_word = 8'hE1;
		16'h51BE: out_word = 8'hCD;
		16'h51BF: out_word = 8'h0C;
		16'h51C0: out_word = 8'h05;
		16'h51C1: out_word = 8'h7E;
		16'h51C2: out_word = 8'hB7;
		16'h51C3: out_word = 8'hCA;
		16'h51C4: out_word = 8'hD3;
		16'h51C5: out_word = 8'h01;
		16'h51C6: out_word = 8'hFE;
		16'h51C7: out_word = 8'h01;
		16'h51C8: out_word = 8'hCC;
		16'h51C9: out_word = 8'h07;
		16'h51CA: out_word = 8'h05;
		16'h51CB: out_word = 8'hC0;
		16'h51CC: out_word = 8'h18;
		16'h51CD: out_word = 8'hE2;
		16'h51CE: out_word = 8'hCD;
		16'h51CF: out_word = 8'h2B;
		16'h51D0: out_word = 8'h04;
		16'h51D1: out_word = 8'h01;
		16'h51D2: out_word = 8'h02;
		16'h51D3: out_word = 8'h00;
		16'h51D4: out_word = 8'hED;
		16'h51D5: out_word = 8'h43;
		16'h51D6: out_word = 8'hDB;
		16'h51D7: out_word = 8'h5C;
		16'h51D8: out_word = 8'h28;
		16'h51D9: out_word = 8'h2B;
		16'h51DA: out_word = 8'hFE;
		16'h51DB: out_word = 8'h23;
		16'h51DC: out_word = 8'h20;
		16'h51DD: out_word = 8'h1A;
		16'h51DE: out_word = 8'h22;
		16'h51DF: out_word = 8'h5D;
		16'h51E0: out_word = 8'h5C;
		16'h51E1: out_word = 8'hCD;
		16'h51E2: out_word = 8'h0B;
		16'h51E3: out_word = 8'h1E;
		16'h51E4: out_word = 8'hCD;
		16'h51E5: out_word = 8'h8C;
		16'h51E6: out_word = 8'h1D;
		16'h51E7: out_word = 8'hFE;
		16'h51E8: out_word = 8'h0D;
		16'h51E9: out_word = 8'h28;
		16'h51EA: out_word = 8'h1A;
		16'h51EB: out_word = 8'hFE;
		16'h51EC: out_word = 8'h2C;
		16'h51ED: out_word = 8'hC2;
		16'h51EE: out_word = 8'h1A;
		16'h51EF: out_word = 8'h1D;
		16'h51F0: out_word = 8'hCD;
		16'h51F1: out_word = 8'h2A;
		16'h51F2: out_word = 8'h1E;
		16'h51F3: out_word = 8'hCD;
		16'h51F4: out_word = 8'hBD;
		16'h51F5: out_word = 8'h1D;
		16'h51F6: out_word = 8'h18;
		16'h51F7: out_word = 8'h03;
		16'h51F8: out_word = 8'hCD;
		16'h51F9: out_word = 8'hDF;
		16'h51FA: out_word = 8'h1D;
		16'h51FB: out_word = 8'hCD;
		16'h51FC: out_word = 8'h75;
		16'h51FD: out_word = 8'h1D;
		16'h51FE: out_word = 8'hCD;
		16'h51FF: out_word = 8'hB5;
		16'h5200: out_word = 8'h1D;
		16'h5201: out_word = 8'hEB;
		16'h5202: out_word = 8'hCD;
		16'h5203: out_word = 8'h81;
		16'h5204: out_word = 8'h1C;
		16'h5205: out_word = 8'hCD;
		16'h5206: out_word = 8'h75;
		16'h5207: out_word = 8'h1D;
		16'h5208: out_word = 8'h3A;
		16'h5209: out_word = 8'hF6;
		16'h520A: out_word = 8'h5C;
		16'h520B: out_word = 8'h32;
		16'h520C: out_word = 8'hF9;
		16'h520D: out_word = 8'h5C;
		16'h520E: out_word = 8'hCD;
		16'h520F: out_word = 8'h05;
		16'h5210: out_word = 8'h04;
		16'h5211: out_word = 8'h3A;
		16'h5212: out_word = 8'hDB;
		16'h5213: out_word = 8'h5C;
		16'h5214: out_word = 8'hFE;
		16'h5215: out_word = 8'h02;
		16'h5216: out_word = 8'hF5;
		16'h5217: out_word = 8'hCC;
		16'h5218: out_word = 8'h97;
		16'h5219: out_word = 8'h1D;
		16'h521A: out_word = 8'hF1;
		16'h521B: out_word = 8'hFE;
		16'h521C: out_word = 8'h11;
		16'h521D: out_word = 8'hD2;
		16'h521E: out_word = 8'h1A;
		16'h521F: out_word = 8'h1D;
		16'h5220: out_word = 8'hCD;
		16'h5221: out_word = 8'h84;
		16'h5222: out_word = 8'h1D;
		16'h5223: out_word = 8'h3E;
		16'h5224: out_word = 8'hFF;
		16'h5225: out_word = 8'h32;
		16'h5226: out_word = 8'hF8;
		16'h5227: out_word = 8'h5C;
		16'h5228: out_word = 8'hCD;
		16'h5229: out_word = 8'h51;
		16'h522A: out_word = 8'h11;
		16'h522B: out_word = 8'hCD;
		16'h522C: out_word = 8'hF6;
		16'h522D: out_word = 8'h3B;
		16'h522E: out_word = 8'hED;
		16'h522F: out_word = 8'h5B;
		16'h5230: out_word = 8'hCF;
		16'h5231: out_word = 8'h5C;
		16'h5232: out_word = 8'h01;
		16'h5233: out_word = 8'h20;
		16'h5234: out_word = 8'h00;
		16'h5235: out_word = 8'hED;
		16'h5236: out_word = 8'hB0;
		16'h5237: out_word = 8'hCD;
		16'h5238: out_word = 8'hE8;
		16'h5239: out_word = 8'h03;
		16'h523A: out_word = 8'h21;
		16'h523B: out_word = 8'h25;
		16'h523C: out_word = 8'h5D;
		16'h523D: out_word = 8'hE5;
		16'h523E: out_word = 8'h21;
		16'h523F: out_word = 8'hB3;
		16'h5240: out_word = 8'h10;
		16'h5241: out_word = 8'hC5;
		16'h5242: out_word = 8'hDF;
		16'h5243: out_word = 8'h2A;
		16'h5244: out_word = 8'hCF;
		16'h5245: out_word = 8'h5C;
		16'h5246: out_word = 8'h01;
		16'h5247: out_word = 8'h14;
		16'h5248: out_word = 8'h00;
		16'h5249: out_word = 8'h09;
		16'h524A: out_word = 8'hDF;
		16'h524B: out_word = 8'h21;
		16'h524C: out_word = 8'hBA;
		16'h524D: out_word = 8'h10;
		16'h524E: out_word = 8'hDF;
		16'h524F: out_word = 8'h3A;
		16'h5250: out_word = 8'hF6;
		16'h5251: out_word = 8'h5C;
		16'h5252: out_word = 8'hC6;
		16'h5253: out_word = 8'h41;
		16'h5254: out_word = 8'hCD;
		16'h5255: out_word = 8'h82;
		16'h5256: out_word = 8'h3D;
		16'h5257: out_word = 8'hCD;
		16'h5258: out_word = 8'h80;
		16'h5259: out_word = 8'h3D;
		16'h525A: out_word = 8'h2A;
		16'h525B: out_word = 8'hCF;
		16'h525C: out_word = 8'h5C;
		16'h525D: out_word = 8'h01;
		16'h525E: out_word = 8'h03;
		16'h525F: out_word = 8'h00;
		16'h5260: out_word = 8'h09;
		16'h5261: out_word = 8'h7E;
		16'h5262: out_word = 8'h2A;
		16'h5263: out_word = 8'hCF;
		16'h5264: out_word = 8'h5C;
		16'h5265: out_word = 8'h01;
		16'h5266: out_word = 8'h13;
		16'h5267: out_word = 8'h00;
		16'h5268: out_word = 8'h09;
		16'h5269: out_word = 8'h96;
		16'h526A: out_word = 8'hE5;
		16'h526B: out_word = 8'hCD;
		16'h526C: out_word = 8'hA3;
		16'h526D: out_word = 8'h1D;
		16'h526E: out_word = 8'h21;
		16'h526F: out_word = 8'hAA;
		16'h5270: out_word = 8'h10;
		16'h5271: out_word = 8'hDF;
		16'h5272: out_word = 8'h2A;
		16'h5273: out_word = 8'hCF;
		16'h5274: out_word = 8'h5C;
		16'h5275: out_word = 8'h01;
		16'h5276: out_word = 8'h02;
		16'h5277: out_word = 8'h00;
		16'h5278: out_word = 8'h09;
		16'h5279: out_word = 8'h7E;
		16'h527A: out_word = 8'h21;
		16'h527B: out_word = 8'hCE;
		16'h527C: out_word = 8'h10;
		16'h527D: out_word = 8'hFE;
		16'h527E: out_word = 8'h19;
		16'h527F: out_word = 8'h28;
		16'h5280: out_word = 8'h11;
		16'h5281: out_word = 8'h21;
		16'h5282: out_word = 8'hE2;
		16'h5283: out_word = 8'h10;
		16'h5284: out_word = 8'hFE;
		16'h5285: out_word = 8'h18;
		16'h5286: out_word = 8'h28;
		16'h5287: out_word = 8'h0A;
		16'h5288: out_word = 8'h21;
		16'h5289: out_word = 8'hF6;
		16'h528A: out_word = 8'h10;
		16'h528B: out_word = 8'hFE;
		16'h528C: out_word = 8'h17;
		16'h528D: out_word = 8'h28;
		16'h528E: out_word = 8'h03;
		16'h528F: out_word = 8'h21;
		16'h5290: out_word = 8'h0A;
		16'h5291: out_word = 8'h11;
		16'h5292: out_word = 8'hDF;
		16'h5293: out_word = 8'hE1;
		16'h5294: out_word = 8'h4E;
		16'h5295: out_word = 8'hCD;
		16'h5296: out_word = 8'hA4;
		16'h5297: out_word = 8'h1D;
		16'h5298: out_word = 8'h21;
		16'h5299: out_word = 8'hA5;
		16'h529A: out_word = 8'h10;
		16'h529B: out_word = 8'hDF;
		16'h529C: out_word = 8'h21;
		16'h529D: out_word = 8'h1E;
		16'h529E: out_word = 8'h11;
		16'h529F: out_word = 8'hDF;
		16'h52A0: out_word = 8'h2A;
		16'h52A1: out_word = 8'hCF;
		16'h52A2: out_word = 8'h5C;
		16'h52A3: out_word = 8'h01;
		16'h52A4: out_word = 8'h04;
		16'h52A5: out_word = 8'h00;
		16'h52A6: out_word = 8'h09;
		16'h52A7: out_word = 8'h4E;
		16'h52A8: out_word = 8'h23;
		16'h52A9: out_word = 8'h46;
		16'h52AA: out_word = 8'hCD;
		16'h52AB: out_word = 8'hA9;
		16'h52AC: out_word = 8'h1D;
		16'h52AD: out_word = 8'h21;
		16'h52AE: out_word = 8'h2E;
		16'h52AF: out_word = 8'h11;
		16'h52B0: out_word = 8'hDF;
		16'h52B1: out_word = 8'hC1;
		16'h52B2: out_word = 8'hE1;
		16'h52B3: out_word = 8'h06;
		16'h52B4: out_word = 8'h10;
		16'h52B5: out_word = 8'hCD;
		16'h52B6: out_word = 8'hB0;
		16'h52B7: out_word = 8'h11;
		16'h52B8: out_word = 8'hCD;
		16'h52B9: out_word = 8'h80;
		16'h52BA: out_word = 8'h3D;
		16'h52BB: out_word = 8'hC5;
		16'h52BC: out_word = 8'hE5;
		16'h52BD: out_word = 8'hCD;
		16'h52BE: out_word = 8'h38;
		16'h52BF: out_word = 8'h29;
		16'h52C0: out_word = 8'h01;
		16'h52C1: out_word = 8'h0D;
		16'h52C2: out_word = 8'h00;
		16'h52C3: out_word = 8'hE1;
		16'h52C4: out_word = 8'hE5;
		16'h52C5: out_word = 8'h09;
		16'h52C6: out_word = 8'h4E;
		16'h52C7: out_word = 8'hC5;
		16'h52C8: out_word = 8'h79;
		16'h52C9: out_word = 8'h06;
		16'h52CA: out_word = 8'h02;
		16'h52CB: out_word = 8'hFE;
		16'h52CC: out_word = 8'h0A;
		16'h52CD: out_word = 8'h38;
		16'h52CE: out_word = 8'h01;
		16'h52CF: out_word = 8'h05;
		16'h52D0: out_word = 8'hFE;
		16'h52D1: out_word = 8'h64;
		16'h52D2: out_word = 8'h30;
		16'h52D3: out_word = 8'h05;
		16'h52D4: out_word = 8'h3E;
		16'h52D5: out_word = 8'h20;
		16'h52D6: out_word = 8'hD7;
		16'h52D7: out_word = 8'h10;
		16'h52D8: out_word = 8'hFB;
		16'h52D9: out_word = 8'hC1;
		16'h52DA: out_word = 8'hCD;
		16'h52DB: out_word = 8'hA9;
		16'h52DC: out_word = 8'h1D;
		16'h52DD: out_word = 8'h21;
		16'h52DE: out_word = 8'hCA;
		16'h52DF: out_word = 8'h10;
		16'h52E0: out_word = 8'hDF;
		16'h52E1: out_word = 8'hE1;
		16'h52E2: out_word = 8'hE5;
		16'h52E3: out_word = 8'h01;
		16'h52E4: out_word = 8'h09;
		16'h52E5: out_word = 8'h00;
		16'h52E6: out_word = 8'h09;
		16'h52E7: out_word = 8'h5E;
		16'h52E8: out_word = 8'h23;
		16'h52E9: out_word = 8'h56;
		16'h52EA: out_word = 8'hE5;
		16'h52EB: out_word = 8'hEB;
		16'h52EC: out_word = 8'hCD;
		16'h52ED: out_word = 8'h5D;
		16'h52EE: out_word = 8'h11;
		16'h52EF: out_word = 8'h3E;
		16'h52F0: out_word = 8'h20;
		16'h52F1: out_word = 8'hCD;
		16'h52F2: out_word = 8'h82;
		16'h52F3: out_word = 8'h3D;
		16'h52F4: out_word = 8'hE1;
		16'h52F5: out_word = 8'h23;
		16'h52F6: out_word = 8'h5E;
		16'h52F7: out_word = 8'h23;
		16'h52F8: out_word = 8'h56;
		16'h52F9: out_word = 8'hEB;
		16'h52FA: out_word = 8'hCD;
		16'h52FB: out_word = 8'h5D;
		16'h52FC: out_word = 8'h11;
		16'h52FD: out_word = 8'hE1;
		16'h52FE: out_word = 8'hE5;
		16'h52FF: out_word = 8'h01;
		16'h5300: out_word = 8'h08;
		16'h5301: out_word = 8'h00;
		16'h5302: out_word = 8'h09;
		16'h5303: out_word = 8'h7E;
		16'h5304: out_word = 8'hFE;
		16'h5305: out_word = 8'h42;
		16'h5306: out_word = 8'hCC;
		16'h5307: out_word = 8'h1B;
		16'h5308: out_word = 8'h13;
		16'h5309: out_word = 8'hE1;
		16'h530A: out_word = 8'hC1;
		16'h530B: out_word = 8'h11;
		16'h530C: out_word = 8'h10;
		16'h530D: out_word = 8'h00;
		16'h530E: out_word = 8'h19;
		16'h530F: out_word = 8'h10;
		16'h5310: out_word = 8'hA4;
		16'h5311: out_word = 8'hE5;
		16'h5312: out_word = 8'hCD;
		16'h5313: out_word = 8'h80;
		16'h5314: out_word = 8'h3D;
		16'h5315: out_word = 8'hCD;
		16'h5316: out_word = 8'h80;
		16'h5317: out_word = 8'h3D;
		16'h5318: out_word = 8'hC3;
		16'h5319: out_word = 8'h3E;
		16'h531A: out_word = 8'h12;
		16'h531B: out_word = 8'h01;
		16'h531C: out_word = 8'h05;
		16'h531D: out_word = 8'h00;
		16'h531E: out_word = 8'h09;
		16'h531F: out_word = 8'h46;
		16'h5320: out_word = 8'h23;
		16'h5321: out_word = 8'h5E;
		16'h5322: out_word = 8'h23;
		16'h5323: out_word = 8'h56;
		16'h5324: out_word = 8'h05;
		16'h5325: out_word = 8'h28;
		16'h5326: out_word = 8'h0E;
		16'h5327: out_word = 8'h05;
		16'h5328: out_word = 8'h28;
		16'h5329: out_word = 8'h0B;
		16'h532A: out_word = 8'h3E;
		16'h532B: out_word = 8'h10;
		16'h532C: out_word = 8'h1C;
		16'h532D: out_word = 8'hBB;
		16'h532E: out_word = 8'h20;
		16'h532F: out_word = 8'h03;
		16'h5330: out_word = 8'h1E;
		16'h5331: out_word = 8'h00;
		16'h5332: out_word = 8'h14;
		16'h5333: out_word = 8'h10;
		16'h5334: out_word = 8'hF7;
		16'h5335: out_word = 8'h2A;
		16'h5336: out_word = 8'hCF;
		16'h5337: out_word = 8'h5C;
		16'h5338: out_word = 8'h01;
		16'h5339: out_word = 8'h21;
		16'h533A: out_word = 8'h00;
		16'h533B: out_word = 8'h09;
		16'h533C: out_word = 8'h06;
		16'h533D: out_word = 8'h02;
		16'h533E: out_word = 8'hE5;
		16'h533F: out_word = 8'hCD;
		16'h5340: out_word = 8'h3D;
		16'h5341: out_word = 8'h1E;
		16'h5342: out_word = 8'h3E;
		16'h5343: out_word = 8'h80;
		16'h5344: out_word = 8'hE1;
		16'h5345: out_word = 8'h01;
		16'h5346: out_word = 8'h00;
		16'h5347: out_word = 8'h02;
		16'h5348: out_word = 8'hED;
		16'h5349: out_word = 8'hB1;
		16'h534A: out_word = 8'h7E;
		16'h534B: out_word = 8'hFE;
		16'h534C: out_word = 8'hAA;
		16'h534D: out_word = 8'hC0;
		16'h534E: out_word = 8'h23;
		16'h534F: out_word = 8'h4E;
		16'h5350: out_word = 8'h23;
		16'h5351: out_word = 8'h46;
		16'h5352: out_word = 8'h78;
		16'h5353: out_word = 8'hB1;
		16'h5354: out_word = 8'hC8;
		16'h5355: out_word = 8'hC5;
		16'h5356: out_word = 8'h3E;
		16'h5357: out_word = 8'h20;
		16'h5358: out_word = 8'hCD;
		16'h5359: out_word = 8'h82;
		16'h535A: out_word = 8'h3D;
		16'h535B: out_word = 8'hC1;
		16'h535C: out_word = 8'hCD;
		16'h535D: out_word = 8'hA9;
		16'h535E: out_word = 8'h1D;
		16'h535F: out_word = 8'hC9;
		16'h5360: out_word = 8'hCD;
		16'h5361: out_word = 8'hC5;
		16'h5362: out_word = 8'h1D;
		16'h5363: out_word = 8'hCD;
		16'h5364: out_word = 8'h2A;
		16'h5365: out_word = 8'h1E;
		16'h5366: out_word = 8'hCD;
		16'h5367: out_word = 8'hBD;
		16'h5368: out_word = 8'h1D;
		16'h5369: out_word = 8'hCD;
		16'h536A: out_word = 8'h75;
		16'h536B: out_word = 8'h1D;
		16'h536C: out_word = 8'hCD;
		16'h536D: out_word = 8'h6F;
		16'h536E: out_word = 8'h16;
		16'h536F: out_word = 8'h21;
		16'h5370: out_word = 8'hAA;
		16'h5371: out_word = 8'h27;
		16'h5372: out_word = 8'hCD;
		16'h5373: out_word = 8'h07;
		16'h5374: out_word = 8'h27;
		16'h5375: out_word = 8'hCD;
		16'h5376: out_word = 8'h52;
		16'h5377: out_word = 8'h10;
		16'h5378: out_word = 8'hFE;
		16'h5379: out_word = 8'h59;
		16'h537A: out_word = 8'h20;
		16'h537B: out_word = 8'hF9;
		16'h537C: out_word = 8'hCD;
		16'h537D: out_word = 8'h9F;
		16'h537E: out_word = 8'h1D;
		16'h537F: out_word = 8'hCD;
		16'h5380: out_word = 8'h2E;
		16'h5381: out_word = 8'h10;
		16'h5382: out_word = 8'hCD;
		16'h5383: out_word = 8'hB0;
		16'h5384: out_word = 8'h1C;
		16'h5385: out_word = 8'hC2;
		16'h5386: out_word = 8'hD9;
		16'h5387: out_word = 8'h03;
		16'h5388: out_word = 8'hCD;
		16'h5389: out_word = 8'hB7;
		16'h538A: out_word = 8'h13;
		16'h538B: out_word = 8'h3A;
		16'h538C: out_word = 8'hE5;
		16'h538D: out_word = 8'h5C;
		16'h538E: out_word = 8'hFE;
		16'h538F: out_word = 8'h23;
		16'h5390: out_word = 8'hC2;
		16'h5391: out_word = 8'hE1;
		16'h5392: out_word = 8'h03;
		16'h5393: out_word = 8'h3E;
		16'h5394: out_word = 8'h0A;
		16'h5395: out_word = 8'h32;
		16'h5396: out_word = 8'h06;
		16'h5397: out_word = 8'h5D;
		16'h5398: out_word = 8'h21;
		16'h5399: out_word = 8'hE6;
		16'h539A: out_word = 8'h5C;
		16'h539B: out_word = 8'h34;
		16'h539C: out_word = 8'hCD;
		16'h539D: out_word = 8'h97;
		16'h539E: out_word = 8'h1D;
		16'h539F: out_word = 8'h21;
		16'h53A0: out_word = 8'hAA;
		16'h53A1: out_word = 8'h27;
		16'h53A2: out_word = 8'hCD;
		16'h53A3: out_word = 8'h07;
		16'h53A4: out_word = 8'h27;
		16'h53A5: out_word = 8'hCD;
		16'h53A6: out_word = 8'h52;
		16'h53A7: out_word = 8'h10;
		16'h53A8: out_word = 8'hFE;
		16'h53A9: out_word = 8'h59;
		16'h53AA: out_word = 8'h20;
		16'h53AB: out_word = 8'hF9;
		16'h53AC: out_word = 8'hCD;
		16'h53AD: out_word = 8'hB3;
		16'h53AE: out_word = 8'h1C;
		16'h53AF: out_word = 8'hC2;
		16'h53B0: out_word = 8'hE1;
		16'h53B1: out_word = 8'h03;
		16'h53B2: out_word = 8'hCD;
		16'h53B3: out_word = 8'hB7;
		16'h53B4: out_word = 8'h13;
		16'h53B5: out_word = 8'h18;
		16'h53B6: out_word = 8'hDC;
		16'h53B7: out_word = 8'hCD;
		16'h53B8: out_word = 8'h5D;
		16'h53B9: out_word = 8'h16;
		16'h53BA: out_word = 8'h21;
		16'h53BB: out_word = 8'hE6;
		16'h53BC: out_word = 8'h5C;
		16'h53BD: out_word = 8'h11;
		16'h53BE: out_word = 8'hED;
		16'h53BF: out_word = 8'h5C;
		16'h53C0: out_word = 8'h01;
		16'h53C1: out_word = 8'h07;
		16'h53C2: out_word = 8'h00;
		16'h53C3: out_word = 8'hED;
		16'h53C4: out_word = 8'hB0;
		16'h53C5: out_word = 8'h3A;
		16'h53C6: out_word = 8'hF1;
		16'h53C7: out_word = 8'h5C;
		16'h53C8: out_word = 8'h32;
		16'h53C9: out_word = 8'h10;
		16'h53CA: out_word = 8'h5D;
		16'h53CB: out_word = 8'hCD;
		16'h53CC: out_word = 8'h05;
		16'h53CD: out_word = 8'h04;
		16'h53CE: out_word = 8'hCD;
		16'h53CF: out_word = 8'h11;
		16'h53D0: out_word = 8'h3E;
		16'h53D1: out_word = 8'h32;
		16'h53D2: out_word = 8'hD9;
		16'h53D3: out_word = 8'h5C;
		16'h53D4: out_word = 8'h3E;
		16'h53D5: out_word = 8'hFF;
		16'h53D6: out_word = 8'h32;
		16'h53D7: out_word = 8'h21;
		16'h53D8: out_word = 8'h5D;
		16'h53D9: out_word = 8'hCD;
		16'h53DA: out_word = 8'h51;
		16'h53DB: out_word = 8'h14;
		16'h53DC: out_word = 8'h2A;
		16'h53DD: out_word = 8'h1F;
		16'h53DE: out_word = 8'h5D;
		16'h53DF: out_word = 8'h22;
		16'h53E0: out_word = 8'hEB;
		16'h53E1: out_word = 8'h5C;
		16'h53E2: out_word = 8'h2A;
		16'h53E3: out_word = 8'hF4;
		16'h53E4: out_word = 8'h5C;
		16'h53E5: out_word = 8'h22;
		16'h53E6: out_word = 8'h06;
		16'h53E7: out_word = 8'h5E;
		16'h53E8: out_word = 8'h21;
		16'h53E9: out_word = 8'h09;
		16'h53EA: out_word = 8'h5E;
		16'h53EB: out_word = 8'h34;
		16'h53EC: out_word = 8'h4E;
		16'h53ED: out_word = 8'h0D;
		16'h53EE: out_word = 8'h06;
		16'h53EF: out_word = 8'h00;
		16'h53F0: out_word = 8'hC5;
		16'h53F1: out_word = 8'h11;
		16'h53F2: out_word = 8'h09;
		16'h53F3: out_word = 8'h00;
		16'h53F4: out_word = 8'hED;
		16'h53F5: out_word = 8'h53;
		16'h53F6: out_word = 8'hF4;
		16'h53F7: out_word = 8'h5C;
		16'h53F8: out_word = 8'hCD;
		16'h53F9: out_word = 8'h43;
		16'h53FA: out_word = 8'h1E;
		16'h53FB: out_word = 8'hC1;
		16'h53FC: out_word = 8'hCD;
		16'h53FD: out_word = 8'h6B;
		16'h53FE: out_word = 8'h16;
		16'h53FF: out_word = 8'hCD;
		16'h5400: out_word = 8'h43;
		16'h5401: out_word = 8'h1E;
		16'h5402: out_word = 8'hC9;
		16'h5403: out_word = 8'hAF;
		16'h5404: out_word = 8'h32;
		16'h5405: out_word = 8'h21;
		16'h5406: out_word = 8'h5D;
		16'h5407: out_word = 8'hCD;
		16'h5408: out_word = 8'h05;
		16'h5409: out_word = 8'h04;
		16'h540A: out_word = 8'hCD;
		16'h540B: out_word = 8'h11;
		16'h540C: out_word = 8'h3E;
		16'h540D: out_word = 8'h32;
		16'h540E: out_word = 8'hDA;
		16'h540F: out_word = 8'h5C;
		16'h5410: out_word = 8'hCD;
		16'h5411: out_word = 8'hB3;
		16'h5412: out_word = 8'h1C;
		16'h5413: out_word = 8'hCA;
		16'h5414: out_word = 8'h50;
		16'h5415: out_word = 8'h1C;
		16'h5416: out_word = 8'hCD;
		16'h5417: out_word = 8'hFD;
		16'h5418: out_word = 8'h03;
		16'h5419: out_word = 8'h3A;
		16'h541A: out_word = 8'h09;
		16'h541B: out_word = 8'h5E;
		16'h541C: out_word = 8'hFE;
		16'h541D: out_word = 8'h80;
		16'h541E: out_word = 8'hCA;
		16'h541F: out_word = 8'h23;
		16'h5420: out_word = 8'h27;
		16'h5421: out_word = 8'h21;
		16'h5422: out_word = 8'hED;
		16'h5423: out_word = 8'h5C;
		16'h5424: out_word = 8'h11;
		16'h5425: out_word = 8'hE6;
		16'h5426: out_word = 8'h5C;
		16'h5427: out_word = 8'h01;
		16'h5428: out_word = 8'h07;
		16'h5429: out_word = 8'h00;
		16'h542A: out_word = 8'hED;
		16'h542B: out_word = 8'hB0;
		16'h542C: out_word = 8'hCD;
		16'h542D: out_word = 8'hFD;
		16'h542E: out_word = 8'h03;
		16'h542F: out_word = 8'h3A;
		16'h5430: out_word = 8'h10;
		16'h5431: out_word = 8'h5D;
		16'h5432: out_word = 8'h32;
		16'h5433: out_word = 8'hEA;
		16'h5434: out_word = 8'h5C;
		16'h5435: out_word = 8'hED;
		16'h5436: out_word = 8'h5B;
		16'h5437: out_word = 8'hEA;
		16'h5438: out_word = 8'h5C;
		16'h5439: out_word = 8'h16;
		16'h543A: out_word = 8'h00;
		16'h543B: out_word = 8'hB7;
		16'h543C: out_word = 8'h2A;
		16'h543D: out_word = 8'h0A;
		16'h543E: out_word = 8'h5E;
		16'h543F: out_word = 8'hED;
		16'h5440: out_word = 8'h52;
		16'h5441: out_word = 8'hDA;
		16'h5442: out_word = 8'h45;
		16'h5443: out_word = 8'h1C;
		16'h5444: out_word = 8'h22;
		16'h5445: out_word = 8'h0A;
		16'h5446: out_word = 8'h5E;
		16'h5447: out_word = 8'h2A;
		16'h5448: out_word = 8'h06;
		16'h5449: out_word = 8'h5E;
		16'h544A: out_word = 8'h22;
		16'h544B: out_word = 8'hEB;
		16'h544C: out_word = 8'h5C;
		16'h544D: out_word = 8'h22;
		16'h544E: out_word = 8'h1F;
		16'h544F: out_word = 8'h5D;
		16'h5450: out_word = 8'hC9;
		16'h5451: out_word = 8'h3A;
		16'h5452: out_word = 8'hF1;
		16'h5453: out_word = 8'h5C;
		16'h5454: out_word = 8'hB7;
		16'h5455: out_word = 8'hC8;
		16'h5456: out_word = 8'h3A;
		16'h5457: out_word = 8'h21;
		16'h5458: out_word = 8'h5D;
		16'h5459: out_word = 8'hB7;
		16'h545A: out_word = 8'h20;
		16'h545B: out_word = 8'h13;
		16'h545C: out_word = 8'hCD;
		16'h545D: out_word = 8'h97;
		16'h545E: out_word = 8'h1D;
		16'h545F: out_word = 8'h21;
		16'h5460: out_word = 8'hAA;
		16'h5461: out_word = 8'h27;
		16'h5462: out_word = 8'hCD;
		16'h5463: out_word = 8'h07;
		16'h5464: out_word = 8'h27;
		16'h5465: out_word = 8'hCD;
		16'h5466: out_word = 8'h52;
		16'h5467: out_word = 8'h10;
		16'h5468: out_word = 8'hFE;
		16'h5469: out_word = 8'h59;
		16'h546A: out_word = 8'h20;
		16'h546B: out_word = 8'hF9;
		16'h546C: out_word = 8'hCD;
		16'h546D: out_word = 8'h9F;
		16'h546E: out_word = 8'h1D;
		16'h546F: out_word = 8'h3A;
		16'h5470: out_word = 8'hF1;
		16'h5471: out_word = 8'h5C;
		16'h5472: out_word = 8'hB7;
		16'h5473: out_word = 8'hC8;
		16'h5474: out_word = 8'hE5;
		16'h5475: out_word = 8'h21;
		16'h5476: out_word = 8'h23;
		16'h5477: out_word = 8'h5D;
		16'h5478: out_word = 8'h96;
		16'h5479: out_word = 8'hE1;
		16'h547A: out_word = 8'h30;
		16'h547B: out_word = 8'h4F;
		16'h547C: out_word = 8'h3A;
		16'h547D: out_word = 8'hF1;
		16'h547E: out_word = 8'h5C;
		16'h547F: out_word = 8'h47;
		16'h5480: out_word = 8'hAF;
		16'h5481: out_word = 8'h32;
		16'h5482: out_word = 8'hF1;
		16'h5483: out_word = 8'h5C;
		16'h5484: out_word = 8'hC5;
		16'h5485: out_word = 8'h32;
		16'h5486: out_word = 8'hCE;
		16'h5487: out_word = 8'h5C;
		16'h5488: out_word = 8'h2A;
		16'h5489: out_word = 8'hCF;
		16'h548A: out_word = 8'h5C;
		16'h548B: out_word = 8'hE5;
		16'h548C: out_word = 8'hED;
		16'h548D: out_word = 8'h5B;
		16'h548E: out_word = 8'hF2;
		16'h548F: out_word = 8'h5C;
		16'h5490: out_word = 8'hCD;
		16'h5491: out_word = 8'hD8;
		16'h5492: out_word = 8'h14;
		16'h5493: out_word = 8'hCD;
		16'h5494: out_word = 8'h3D;
		16'h5495: out_word = 8'h1E;
		16'h5496: out_word = 8'h2A;
		16'h5497: out_word = 8'hF4;
		16'h5498: out_word = 8'h5C;
		16'h5499: out_word = 8'h22;
		16'h549A: out_word = 8'hF2;
		16'h549B: out_word = 8'h5C;
		16'h549C: out_word = 8'hCD;
		16'h549D: out_word = 8'h97;
		16'h549E: out_word = 8'h1D;
		16'h549F: out_word = 8'h21;
		16'h54A0: out_word = 8'h85;
		16'h54A1: out_word = 8'h27;
		16'h54A2: out_word = 8'hCD;
		16'h54A3: out_word = 8'h07;
		16'h54A4: out_word = 8'h27;
		16'h54A5: out_word = 8'hCD;
		16'h54A6: out_word = 8'h52;
		16'h54A7: out_word = 8'h10;
		16'h54A8: out_word = 8'hFE;
		16'h54A9: out_word = 8'h59;
		16'h54AA: out_word = 8'h20;
		16'h54AB: out_word = 8'hF9;
		16'h54AC: out_word = 8'hCD;
		16'h54AD: out_word = 8'h9F;
		16'h54AE: out_word = 8'h1D;
		16'h54AF: out_word = 8'h3A;
		16'h54B0: out_word = 8'h21;
		16'h54B1: out_word = 8'h5D;
		16'h54B2: out_word = 8'hB7;
		16'h54B3: out_word = 8'hC4;
		16'h54B4: out_word = 8'h03;
		16'h54B5: out_word = 8'h14;
		16'h54B6: out_word = 8'hE1;
		16'h54B7: out_word = 8'hC1;
		16'h54B8: out_word = 8'hED;
		16'h54B9: out_word = 8'h5B;
		16'h54BA: out_word = 8'hEB;
		16'h54BB: out_word = 8'h5C;
		16'h54BC: out_word = 8'hCD;
		16'h54BD: out_word = 8'hE4;
		16'h54BE: out_word = 8'h14;
		16'h54BF: out_word = 8'hCD;
		16'h54C0: out_word = 8'h4D;
		16'h54C1: out_word = 8'h1E;
		16'h54C2: out_word = 8'h2A;
		16'h54C3: out_word = 8'hF4;
		16'h54C4: out_word = 8'h5C;
		16'h54C5: out_word = 8'h22;
		16'h54C6: out_word = 8'hEB;
		16'h54C7: out_word = 8'h5C;
		16'h54C8: out_word = 8'hC3;
		16'h54C9: out_word = 8'h51;
		16'h54CA: out_word = 8'h14;
		16'h54CB: out_word = 8'h32;
		16'h54CC: out_word = 8'hF1;
		16'h54CD: out_word = 8'h5C;
		16'h54CE: out_word = 8'hE5;
		16'h54CF: out_word = 8'h21;
		16'h54D0: out_word = 8'h23;
		16'h54D1: out_word = 8'h5D;
		16'h54D2: out_word = 8'h46;
		16'h54D3: out_word = 8'hE1;
		16'h54D4: out_word = 8'hAF;
		16'h54D5: out_word = 8'hC3;
		16'h54D6: out_word = 8'h84;
		16'h54D7: out_word = 8'h14;
		16'h54D8: out_word = 8'hE5;
		16'h54D9: out_word = 8'hD5;
		16'h54DA: out_word = 8'hCD;
		16'h54DB: out_word = 8'h11;
		16'h54DC: out_word = 8'h3E;
		16'h54DD: out_word = 8'h3A;
		16'h54DE: out_word = 8'hD9;
		16'h54DF: out_word = 8'h5C;
		16'h54E0: out_word = 8'h77;
		16'h54E1: out_word = 8'hD1;
		16'h54E2: out_word = 8'hE1;
		16'h54E3: out_word = 8'hC9;
		16'h54E4: out_word = 8'hE5;
		16'h54E5: out_word = 8'hD5;
		16'h54E6: out_word = 8'hCD;
		16'h54E7: out_word = 8'h11;
		16'h54E8: out_word = 8'h3E;
		16'h54E9: out_word = 8'h3A;
		16'h54EA: out_word = 8'hDA;
		16'h54EB: out_word = 8'h5C;
		16'h54EC: out_word = 8'h77;
		16'h54ED: out_word = 8'hD1;
		16'h54EE: out_word = 8'hE1;
		16'h54EF: out_word = 8'hC9;
		16'h54F0: out_word = 8'hAF;
		16'h54F1: out_word = 8'h32;
		16'h54F2: out_word = 8'h21;
		16'h54F3: out_word = 8'h5D;
		16'h54F4: out_word = 8'hCD;
		16'h54F5: out_word = 8'h05;
		16'h54F6: out_word = 8'h04;
		16'h54F7: out_word = 8'hCD;
		16'h54F8: out_word = 8'h11;
		16'h54F9: out_word = 8'h3E;
		16'h54FA: out_word = 8'h32;
		16'h54FB: out_word = 8'hDA;
		16'h54FC: out_word = 8'h5C;
		16'h54FD: out_word = 8'h3A;
		16'h54FE: out_word = 8'h08;
		16'h54FF: out_word = 8'h5E;
		16'h5500: out_word = 8'h32;
		16'h5501: out_word = 8'hE7;
		16'h5502: out_word = 8'h5C;
		16'h5503: out_word = 8'h21;
		16'h5504: out_word = 8'h80;
		16'h5505: out_word = 8'h02;
		16'h5506: out_word = 8'hFE;
		16'h5507: out_word = 8'h19;
		16'h5508: out_word = 8'h28;
		16'h5509: out_word = 8'h15;
		16'h550A: out_word = 8'h21;
		16'h550B: out_word = 8'h00;
		16'h550C: out_word = 8'h05;
		16'h550D: out_word = 8'hFE;
		16'h550E: out_word = 8'h18;
		16'h550F: out_word = 8'h28;
		16'h5510: out_word = 8'h0E;
		16'h5511: out_word = 8'hFE;
		16'h5512: out_word = 8'h17;
		16'h5513: out_word = 8'h28;
		16'h5514: out_word = 8'h0A;
		16'h5515: out_word = 8'h21;
		16'h5516: out_word = 8'h00;
		16'h5517: out_word = 8'h0A;
		16'h5518: out_word = 8'hFE;
		16'h5519: out_word = 8'h16;
		16'h551A: out_word = 8'h28;
		16'h551B: out_word = 8'h03;
		16'h551C: out_word = 8'hC3;
		16'h551D: out_word = 8'h1A;
		16'h551E: out_word = 8'h1D;
		16'h551F: out_word = 8'h22;
		16'h5520: out_word = 8'hDD;
		16'h5521: out_word = 8'h5C;
		16'h5522: out_word = 8'hED;
		16'h5523: out_word = 8'h4B;
		16'h5524: out_word = 8'hDF;
		16'h5525: out_word = 8'h5C;
		16'h5526: out_word = 8'hED;
		16'h5527: out_word = 8'h42;
		16'h5528: out_word = 8'hDA;
		16'h5529: out_word = 8'h45;
		16'h552A: out_word = 8'h1C;
		16'h552B: out_word = 8'hC9;
		16'h552C: out_word = 8'hCD;
		16'h552D: out_word = 8'h75;
		16'h552E: out_word = 8'h1D;
		16'h552F: out_word = 8'hCD;
		16'h5530: out_word = 8'h6F;
		16'h5531: out_word = 8'h16;
		16'h5532: out_word = 8'h21;
		16'h5533: out_word = 8'h79;
		16'h5534: out_word = 8'h27;
		16'h5535: out_word = 8'hCD;
		16'h5536: out_word = 8'h07;
		16'h5537: out_word = 8'h27;
		16'h5538: out_word = 8'h21;
		16'h5539: out_word = 8'hAA;
		16'h553A: out_word = 8'h27;
		16'h553B: out_word = 8'hCD;
		16'h553C: out_word = 8'h07;
		16'h553D: out_word = 8'h27;
		16'h553E: out_word = 8'hCD;
		16'h553F: out_word = 8'h52;
		16'h5540: out_word = 8'h10;
		16'h5541: out_word = 8'hFE;
		16'h5542: out_word = 8'h59;
		16'h5543: out_word = 8'h20;
		16'h5544: out_word = 8'hF9;
		16'h5545: out_word = 8'hCD;
		16'h5546: out_word = 8'h9F;
		16'h5547: out_word = 8'h1D;
		16'h5548: out_word = 8'h3E;
		16'h5549: out_word = 8'hFF;
		16'h554A: out_word = 8'h32;
		16'h554B: out_word = 8'h21;
		16'h554C: out_word = 8'h5D;
		16'h554D: out_word = 8'hCD;
		16'h554E: out_word = 8'h05;
		16'h554F: out_word = 8'h04;
		16'h5550: out_word = 8'hCD;
		16'h5551: out_word = 8'h11;
		16'h5552: out_word = 8'h3E;
		16'h5553: out_word = 8'h32;
		16'h5554: out_word = 8'hD9;
		16'h5555: out_word = 8'h5C;
		16'h5556: out_word = 8'h3A;
		16'h5557: out_word = 8'h08;
		16'h5558: out_word = 8'h5E;
		16'h5559: out_word = 8'hFE;
		16'h555A: out_word = 8'h19;
		16'h555B: out_word = 8'h21;
		16'h555C: out_word = 8'h80;
		16'h555D: out_word = 8'h02;
		16'h555E: out_word = 8'h28;
		16'h555F: out_word = 8'h15;
		16'h5560: out_word = 8'h21;
		16'h5561: out_word = 8'h00;
		16'h5562: out_word = 8'h05;
		16'h5563: out_word = 8'hFE;
		16'h5564: out_word = 8'h18;
		16'h5565: out_word = 8'h28;
		16'h5566: out_word = 8'h0E;
		16'h5567: out_word = 8'hFE;
		16'h5568: out_word = 8'h17;
		16'h5569: out_word = 8'h28;
		16'h556A: out_word = 8'h0A;
		16'h556B: out_word = 8'h21;
		16'h556C: out_word = 8'h00;
		16'h556D: out_word = 8'h0A;
		16'h556E: out_word = 8'hFE;
		16'h556F: out_word = 8'h16;
		16'h5570: out_word = 8'h28;
		16'h5571: out_word = 8'h03;
		16'h5572: out_word = 8'hC3;
		16'h5573: out_word = 8'h0F;
		16'h5574: out_word = 8'h04;
		16'h5575: out_word = 8'hED;
		16'h5576: out_word = 8'h4B;
		16'h5577: out_word = 8'h0A;
		16'h5578: out_word = 8'h5E;
		16'h5579: out_word = 8'hED;
		16'h557A: out_word = 8'h42;
		16'h557B: out_word = 8'h22;
		16'h557C: out_word = 8'hE5;
		16'h557D: out_word = 8'h5C;
		16'h557E: out_word = 8'h22;
		16'h557F: out_word = 8'hDF;
		16'h5580: out_word = 8'h5C;
		16'h5581: out_word = 8'h21;
		16'h5582: out_word = 8'h00;
		16'h5583: out_word = 8'h00;
		16'h5584: out_word = 8'h22;
		16'h5585: out_word = 8'hE1;
		16'h5586: out_word = 8'h5C;
		16'h5587: out_word = 8'h22;
		16'h5588: out_word = 8'hE3;
		16'h5589: out_word = 8'h5C;
		16'h558A: out_word = 8'hCD;
		16'h558B: out_word = 8'hB8;
		16'h558C: out_word = 8'h15;
		16'h558D: out_word = 8'hCD;
		16'h558E: out_word = 8'h05;
		16'h558F: out_word = 8'h04;
		16'h5590: out_word = 8'h3A;
		16'h5591: out_word = 8'hE7;
		16'h5592: out_word = 8'h5C;
		16'h5593: out_word = 8'h32;
		16'h5594: out_word = 8'h08;
		16'h5595: out_word = 8'h5E;
		16'h5596: out_word = 8'h2A;
		16'h5597: out_word = 8'hDD;
		16'h5598: out_word = 8'h5C;
		16'h5599: out_word = 8'hED;
		16'h559A: out_word = 8'h4B;
		16'h559B: out_word = 8'hDF;
		16'h559C: out_word = 8'h5C;
		16'h559D: out_word = 8'hED;
		16'h559E: out_word = 8'h42;
		16'h559F: out_word = 8'h22;
		16'h55A0: out_word = 8'h0A;
		16'h55A1: out_word = 8'h5E;
		16'h55A2: out_word = 8'hCD;
		16'h55A3: out_word = 8'hE4;
		16'h55A4: out_word = 8'h14;
		16'h55A5: out_word = 8'h11;
		16'h55A6: out_word = 8'h09;
		16'h55A7: out_word = 8'h00;
		16'h55A8: out_word = 8'hED;
		16'h55A9: out_word = 8'h53;
		16'h55AA: out_word = 8'hF4;
		16'h55AB: out_word = 8'h5C;
		16'h55AC: out_word = 8'hCD;
		16'h55AD: out_word = 8'h43;
		16'h55AE: out_word = 8'h1E;
		16'h55AF: out_word = 8'hC3;
		16'h55B0: out_word = 8'hE1;
		16'h55B1: out_word = 8'h03;
		16'h55B2: out_word = 8'h2A;
		16'h55B3: out_word = 8'hE5;
		16'h55B4: out_word = 8'h5C;
		16'h55B5: out_word = 8'h7C;
		16'h55B6: out_word = 8'hB5;
		16'h55B7: out_word = 8'hC9;
		16'h55B8: out_word = 8'hCD;
		16'h55B9: out_word = 8'hB2;
		16'h55BA: out_word = 8'h15;
		16'h55BB: out_word = 8'hC8;
		16'h55BC: out_word = 8'h3A;
		16'h55BD: out_word = 8'h21;
		16'h55BE: out_word = 8'h5D;
		16'h55BF: out_word = 8'hB7;
		16'h55C0: out_word = 8'h20;
		16'h55C1: out_word = 8'h19;
		16'h55C2: out_word = 8'hCD;
		16'h55C3: out_word = 8'h97;
		16'h55C4: out_word = 8'h1D;
		16'h55C5: out_word = 8'h21;
		16'h55C6: out_word = 8'h79;
		16'h55C7: out_word = 8'h27;
		16'h55C8: out_word = 8'hCD;
		16'h55C9: out_word = 8'h07;
		16'h55CA: out_word = 8'h27;
		16'h55CB: out_word = 8'h21;
		16'h55CC: out_word = 8'hAA;
		16'h55CD: out_word = 8'h27;
		16'h55CE: out_word = 8'hCD;
		16'h55CF: out_word = 8'h07;
		16'h55D0: out_word = 8'h27;
		16'h55D1: out_word = 8'hCD;
		16'h55D2: out_word = 8'h52;
		16'h55D3: out_word = 8'h10;
		16'h55D4: out_word = 8'hFE;
		16'h55D5: out_word = 8'h59;
		16'h55D6: out_word = 8'h20;
		16'h55D7: out_word = 8'hF9;
		16'h55D8: out_word = 8'hCD;
		16'h55D9: out_word = 8'h9F;
		16'h55DA: out_word = 8'h1D;
		16'h55DB: out_word = 8'hCD;
		16'h55DC: out_word = 8'hB2;
		16'h55DD: out_word = 8'h15;
		16'h55DE: out_word = 8'hC8;
		16'h55DF: out_word = 8'hC5;
		16'h55E0: out_word = 8'hE5;
		16'h55E1: out_word = 8'h21;
		16'h55E2: out_word = 8'h23;
		16'h55E3: out_word = 8'h5D;
		16'h55E4: out_word = 8'h4E;
		16'h55E5: out_word = 8'h06;
		16'h55E6: out_word = 8'h00;
		16'h55E7: out_word = 8'hE1;
		16'h55E8: out_word = 8'hED;
		16'h55E9: out_word = 8'h42;
		16'h55EA: out_word = 8'hC1;
		16'h55EB: out_word = 8'hD2;
		16'h55EC: out_word = 8'h44;
		16'h55ED: out_word = 8'h16;
		16'h55EE: out_word = 8'hED;
		16'h55EF: out_word = 8'h4B;
		16'h55F0: out_word = 8'hE5;
		16'h55F1: out_word = 8'h5C;
		16'h55F2: out_word = 8'h21;
		16'h55F3: out_word = 8'h00;
		16'h55F4: out_word = 8'h00;
		16'h55F5: out_word = 8'h22;
		16'h55F6: out_word = 8'hE5;
		16'h55F7: out_word = 8'h5C;
		16'h55F8: out_word = 8'hC5;
		16'h55F9: out_word = 8'h2A;
		16'h55FA: out_word = 8'hCF;
		16'h55FB: out_word = 8'h5C;
		16'h55FC: out_word = 8'hE5;
		16'h55FD: out_word = 8'hCD;
		16'h55FE: out_word = 8'hD8;
		16'h55FF: out_word = 8'h14;
		16'h5600: out_word = 8'hED;
		16'h5601: out_word = 8'h5B;
		16'h5602: out_word = 8'hE1;
		16'h5603: out_word = 8'h5C;
		16'h5604: out_word = 8'h41;
		16'h5605: out_word = 8'hCD;
		16'h5606: out_word = 8'h3D;
		16'h5607: out_word = 8'h1E;
		16'h5608: out_word = 8'h2A;
		16'h5609: out_word = 8'hF4;
		16'h560A: out_word = 8'h5C;
		16'h560B: out_word = 8'h22;
		16'h560C: out_word = 8'hE1;
		16'h560D: out_word = 8'h5C;
		16'h560E: out_word = 8'hCD;
		16'h560F: out_word = 8'h97;
		16'h5610: out_word = 8'h1D;
		16'h5611: out_word = 8'h21;
		16'h5612: out_word = 8'h79;
		16'h5613: out_word = 8'h27;
		16'h5614: out_word = 8'hCD;
		16'h5615: out_word = 8'h07;
		16'h5616: out_word = 8'h27;
		16'h5617: out_word = 8'h21;
		16'h5618: out_word = 8'h85;
		16'h5619: out_word = 8'h27;
		16'h561A: out_word = 8'hCD;
		16'h561B: out_word = 8'h07;
		16'h561C: out_word = 8'h27;
		16'h561D: out_word = 8'hCD;
		16'h561E: out_word = 8'h52;
		16'h561F: out_word = 8'h10;
		16'h5620: out_word = 8'hFE;
		16'h5621: out_word = 8'h59;
		16'h5622: out_word = 8'h20;
		16'h5623: out_word = 8'hF9;
		16'h5624: out_word = 8'hCD;
		16'h5625: out_word = 8'h9F;
		16'h5626: out_word = 8'h1D;
		16'h5627: out_word = 8'h3A;
		16'h5628: out_word = 8'h21;
		16'h5629: out_word = 8'h5D;
		16'h562A: out_word = 8'hB7;
		16'h562B: out_word = 8'hC4;
		16'h562C: out_word = 8'hF0;
		16'h562D: out_word = 8'h14;
		16'h562E: out_word = 8'hE1;
		16'h562F: out_word = 8'hC1;
		16'h5630: out_word = 8'hED;
		16'h5631: out_word = 8'h5B;
		16'h5632: out_word = 8'hE3;
		16'h5633: out_word = 8'h5C;
		16'h5634: out_word = 8'h41;
		16'h5635: out_word = 8'hCD;
		16'h5636: out_word = 8'hE4;
		16'h5637: out_word = 8'h14;
		16'h5638: out_word = 8'hCD;
		16'h5639: out_word = 8'h4D;
		16'h563A: out_word = 8'h1E;
		16'h563B: out_word = 8'h2A;
		16'h563C: out_word = 8'hF4;
		16'h563D: out_word = 8'h5C;
		16'h563E: out_word = 8'h22;
		16'h563F: out_word = 8'hE3;
		16'h5640: out_word = 8'h5C;
		16'h5641: out_word = 8'hC3;
		16'h5642: out_word = 8'hB8;
		16'h5643: out_word = 8'h15;
		16'h5644: out_word = 8'h22;
		16'h5645: out_word = 8'hE5;
		16'h5646: out_word = 8'h5C;
		16'h5647: out_word = 8'hE5;
		16'h5648: out_word = 8'h21;
		16'h5649: out_word = 8'h23;
		16'h564A: out_word = 8'h5D;
		16'h564B: out_word = 8'h4E;
		16'h564C: out_word = 8'h06;
		16'h564D: out_word = 8'h00;
		16'h564E: out_word = 8'hE1;
		16'h564F: out_word = 8'hAF;
		16'h5650: out_word = 8'hC3;
		16'h5651: out_word = 8'hF8;
		16'h5652: out_word = 8'h15;
		16'h5653: out_word = 8'hCD;
		16'h5654: out_word = 8'h5D;
		16'h5655: out_word = 8'h16;
		16'h5656: out_word = 8'h3A;
		16'h5657: out_word = 8'hDD;
		16'h5658: out_word = 8'h5C;
		16'h5659: out_word = 8'hFE;
		16'h565A: out_word = 8'h01;
		16'h565B: out_word = 8'hC9;
		16'h565C: out_word = 8'h4F;
		16'h565D: out_word = 8'hAF;
		16'h565E: out_word = 8'hC5;
		16'h565F: out_word = 8'hCD;
		16'h5660: out_word = 8'hE9;
		16'h5661: out_word = 8'h17;
		16'h5662: out_word = 8'hC1;
		16'h5663: out_word = 8'hC9;
		16'h5664: out_word = 8'h4F;
		16'h5665: out_word = 8'hCD;
		16'h5666: out_word = 8'h6B;
		16'h5667: out_word = 8'h16;
		16'h5668: out_word = 8'hC3;
		16'h5669: out_word = 8'h43;
		16'h566A: out_word = 8'h1E;
		16'h566B: out_word = 8'h3E;
		16'h566C: out_word = 8'hFF;
		16'h566D: out_word = 8'h18;
		16'h566E: out_word = 8'hEF;
		16'h566F: out_word = 8'h3E;
		16'h5670: out_word = 8'hFF;
		16'h5671: out_word = 8'h32;
		16'h5672: out_word = 8'h0E;
		16'h5673: out_word = 8'h5D;
		16'h5674: out_word = 8'hCD;
		16'h5675: out_word = 8'h80;
		16'h5676: out_word = 8'h16;
		16'h5677: out_word = 8'h2A;
		16'h5678: out_word = 8'h61;
		16'h5679: out_word = 8'h5C;
		16'h567A: out_word = 8'h22;
		16'h567B: out_word = 8'hCF;
		16'h567C: out_word = 8'h5C;
		16'h567D: out_word = 8'hC3;
		16'h567E: out_word = 8'h23;
		16'h567F: out_word = 8'h1E;
		16'h5680: out_word = 8'hE7;
		16'h5681: out_word = 8'h1A;
		16'h5682: out_word = 8'h1F;
		16'h5683: out_word = 8'h21;
		16'h5684: out_word = 8'hFF;
		16'h5685: out_word = 8'hFF;
		16'h5686: out_word = 8'hED;
		16'h5687: out_word = 8'h42;
		16'h5688: out_word = 8'h7C;
		16'h5689: out_word = 8'hFE;
		16'h568A: out_word = 8'h10;
		16'h568B: out_word = 8'h30;
		16'h568C: out_word = 8'h02;
		16'h568D: out_word = 8'h3E;
		16'h568E: out_word = 8'h11;
		16'h568F: out_word = 8'h3D;
		16'h5690: out_word = 8'h32;
		16'h5691: out_word = 8'h23;
		16'h5692: out_word = 8'h5D;
		16'h5693: out_word = 8'h47;
		16'h5694: out_word = 8'h0E;
		16'h5695: out_word = 8'h00;
		16'h5696: out_word = 8'hC9;
		16'h5697: out_word = 8'h22;
		16'h5698: out_word = 8'hD7;
		16'h5699: out_word = 8'h5C;
		16'h569A: out_word = 8'h22;
		16'h569B: out_word = 8'hDB;
		16'h569C: out_word = 8'h5C;
		16'h569D: out_word = 8'hED;
		16'h569E: out_word = 8'h5B;
		16'h569F: out_word = 8'hEA;
		16'h56A0: out_word = 8'h5C;
		16'h56A1: out_word = 8'h2A;
		16'h56A2: out_word = 8'hD9;
		16'h56A3: out_word = 8'h5C;
		16'h56A4: out_word = 8'h16;
		16'h56A5: out_word = 8'h00;
		16'h56A6: out_word = 8'h19;
		16'h56A7: out_word = 8'h22;
		16'h56A8: out_word = 8'hD9;
		16'h56A9: out_word = 8'h5C;
		16'h56AA: out_word = 8'hC9;
		16'h56AB: out_word = 8'hCD;
		16'h56AC: out_word = 8'h2B;
		16'h56AD: out_word = 8'h04;
		16'h56AE: out_word = 8'hC2;
		16'h56AF: out_word = 8'h75;
		16'h56B0: out_word = 8'h17;
		16'h56B1: out_word = 8'hCD;
		16'h56B2: out_word = 8'h75;
		16'h56B3: out_word = 8'h1D;
		16'h56B4: out_word = 8'hCD;
		16'h56B5: out_word = 8'h6F;
		16'h56B6: out_word = 8'h16;
		16'h56B7: out_word = 8'h2A;
		16'h56B8: out_word = 8'hCF;
		16'h56B9: out_word = 8'h5C;
		16'h56BA: out_word = 8'h22;
		16'h56BB: out_word = 8'hE1;
		16'h56BC: out_word = 8'h5C;
		16'h56BD: out_word = 8'h11;
		16'h56BE: out_word = 8'h00;
		16'h56BF: out_word = 8'h09;
		16'h56C0: out_word = 8'h19;
		16'h56C1: out_word = 8'h22;
		16'h56C2: out_word = 8'hCF;
		16'h56C3: out_word = 8'h5C;
		16'h56C4: out_word = 8'h3A;
		16'h56C5: out_word = 8'h23;
		16'h56C6: out_word = 8'h5D;
		16'h56C7: out_word = 8'hD6;
		16'h56C8: out_word = 8'h09;
		16'h56C9: out_word = 8'h32;
		16'h56CA: out_word = 8'h23;
		16'h56CB: out_word = 8'h5D;
		16'h56CC: out_word = 8'h2A;
		16'h56CD: out_word = 8'hE1;
		16'h56CE: out_word = 8'h5C;
		16'h56CF: out_word = 8'h11;
		16'h56D0: out_word = 8'h00;
		16'h56D1: out_word = 8'h00;
		16'h56D2: out_word = 8'h06;
		16'h56D3: out_word = 8'h09;
		16'h56D4: out_word = 8'hCD;
		16'h56D5: out_word = 8'h3D;
		16'h56D6: out_word = 8'h1E;
		16'h56D7: out_word = 8'h2A;
		16'h56D8: out_word = 8'hE1;
		16'h56D9: out_word = 8'h5C;
		16'h56DA: out_word = 8'h22;
		16'h56DB: out_word = 8'hDF;
		16'h56DC: out_word = 8'h5C;
		16'h56DD: out_word = 8'h21;
		16'h56DE: out_word = 8'h00;
		16'h56DF: out_word = 8'h01;
		16'h56E0: out_word = 8'h22;
		16'h56E1: out_word = 8'hD7;
		16'h56E2: out_word = 8'h5C;
		16'h56E3: out_word = 8'h22;
		16'h56E4: out_word = 8'hDD;
		16'h56E5: out_word = 8'h5C;
		16'h56E6: out_word = 8'hAF;
		16'h56E7: out_word = 8'h22;
		16'h56E8: out_word = 8'hE3;
		16'h56E9: out_word = 8'h5C;
		16'h56EA: out_word = 8'h32;
		16'h56EB: out_word = 8'hE4;
		16'h56EC: out_word = 8'h5C;
		16'h56ED: out_word = 8'hCD;
		16'h56EE: out_word = 8'h00;
		16'h56EF: out_word = 8'h3B;
		16'h56F0: out_word = 8'hED;
		16'h56F1: out_word = 8'h5B;
		16'h56F2: out_word = 8'hE1;
		16'h56F3: out_word = 8'h5C;
		16'h56F4: out_word = 8'h2A;
		16'h56F5: out_word = 8'hDF;
		16'h56F6: out_word = 8'h5C;
		16'h56F7: out_word = 8'hEB;
		16'h56F8: out_word = 8'h01;
		16'h56F9: out_word = 8'h00;
		16'h56FA: out_word = 8'h08;
		16'h56FB: out_word = 8'h09;
		16'h56FC: out_word = 8'hA7;
		16'h56FD: out_word = 8'hED;
		16'h56FE: out_word = 8'h52;
		16'h56FF: out_word = 8'h2B;
		16'h5700: out_word = 8'h4D;
		16'h5701: out_word = 8'h44;
		16'h5702: out_word = 8'hEB;
		16'h5703: out_word = 8'h54;
		16'h5704: out_word = 8'h5D;
		16'h5705: out_word = 8'h13;
		16'h5706: out_word = 8'h36;
		16'h5707: out_word = 8'h00;
		16'h5708: out_word = 8'hED;
		16'h5709: out_word = 8'hB0;
		16'h570A: out_word = 8'h2A;
		16'h570B: out_word = 8'hE1;
		16'h570C: out_word = 8'h5C;
		16'h570D: out_word = 8'h11;
		16'h570E: out_word = 8'hE1;
		16'h570F: out_word = 8'h08;
		16'h5710: out_word = 8'h19;
		16'h5711: out_word = 8'h5E;
		16'h5712: out_word = 8'h23;
		16'h5713: out_word = 8'h56;
		16'h5714: out_word = 8'hED;
		16'h5715: out_word = 8'h4B;
		16'h5716: out_word = 8'hD7;
		16'h5717: out_word = 8'h5C;
		16'h5718: out_word = 8'h70;
		16'h5719: out_word = 8'h2B;
		16'h571A: out_word = 8'h71;
		16'h571B: out_word = 8'h23;
		16'h571C: out_word = 8'h23;
		16'h571D: out_word = 8'h23;
		16'h571E: out_word = 8'h23;
		16'h571F: out_word = 8'h4E;
		16'h5720: out_word = 8'h23;
		16'h5721: out_word = 8'h46;
		16'h5722: out_word = 8'hEB;
		16'h5723: out_word = 8'h7D;
		16'h5724: out_word = 8'hE6;
		16'h5725: out_word = 8'h0F;
		16'h5726: out_word = 8'h6C;
		16'h5727: out_word = 8'h26;
		16'h5728: out_word = 8'h00;
		16'h5729: out_word = 8'h29;
		16'h572A: out_word = 8'h29;
		16'h572B: out_word = 8'h29;
		16'h572C: out_word = 8'h29;
		16'h572D: out_word = 8'h85;
		16'h572E: out_word = 8'h6F;
		16'h572F: out_word = 8'h09;
		16'h5730: out_word = 8'hED;
		16'h5731: out_word = 8'h4B;
		16'h5732: out_word = 8'hD7;
		16'h5733: out_word = 8'h5C;
		16'h5734: out_word = 8'h22;
		16'h5735: out_word = 8'hD7;
		16'h5736: out_word = 8'h5C;
		16'h5737: out_word = 8'h68;
		16'h5738: out_word = 8'h26;
		16'h5739: out_word = 8'h00;
		16'h573A: out_word = 8'h29;
		16'h573B: out_word = 8'h29;
		16'h573C: out_word = 8'h29;
		16'h573D: out_word = 8'h29;
		16'h573E: out_word = 8'h79;
		16'h573F: out_word = 8'hE6;
		16'h5740: out_word = 8'h0F;
		16'h5741: out_word = 8'h85;
		16'h5742: out_word = 8'h4F;
		16'h5743: out_word = 8'h44;
		16'h5744: out_word = 8'h2A;
		16'h5745: out_word = 8'hD7;
		16'h5746: out_word = 8'h5C;
		16'h5747: out_word = 8'hA7;
		16'h5748: out_word = 8'hED;
		16'h5749: out_word = 8'h42;
		16'h574A: out_word = 8'hEB;
		16'h574B: out_word = 8'h72;
		16'h574C: out_word = 8'h2B;
		16'h574D: out_word = 8'h73;
		16'h574E: out_word = 8'h2B;
		16'h574F: out_word = 8'h3A;
		16'h5750: out_word = 8'hE3;
		16'h5751: out_word = 8'h5C;
		16'h5752: out_word = 8'h77;
		16'h5753: out_word = 8'h11;
		16'h5754: out_word = 8'h10;
		16'h5755: out_word = 8'h00;
		16'h5756: out_word = 8'h19;
		16'h5757: out_word = 8'h36;
		16'h5758: out_word = 8'h00;
		16'h5759: out_word = 8'h2A;
		16'h575A: out_word = 8'hE1;
		16'h575B: out_word = 8'h5C;
		16'h575C: out_word = 8'h11;
		16'h575D: out_word = 8'h00;
		16'h575E: out_word = 8'h00;
		16'h575F: out_word = 8'h06;
		16'h5760: out_word = 8'h09;
		16'h5761: out_word = 8'hCD;
		16'h5762: out_word = 8'h4D;
		16'h5763: out_word = 8'h1E;
		16'h5764: out_word = 8'h3A;
		16'h5765: out_word = 8'h23;
		16'h5766: out_word = 8'h5D;
		16'h5767: out_word = 8'hC6;
		16'h5768: out_word = 8'h09;
		16'h5769: out_word = 8'h47;
		16'h576A: out_word = 8'h0E;
		16'h576B: out_word = 8'h00;
		16'h576C: out_word = 8'h2A;
		16'h576D: out_word = 8'hCF;
		16'h576E: out_word = 8'h5C;
		16'h576F: out_word = 8'hCD;
		16'h5770: out_word = 8'h2E;
		16'h5771: out_word = 8'h1E;
		16'h5772: out_word = 8'hC3;
		16'h5773: out_word = 8'hE1;
		16'h5774: out_word = 8'h03;
		16'h5775: out_word = 8'hCD;
		16'h5776: out_word = 8'hDF;
		16'h5777: out_word = 8'h1D;
		16'h5778: out_word = 8'hCD;
		16'h5779: out_word = 8'h75;
		16'h577A: out_word = 8'h1D;
		16'h577B: out_word = 8'hCD;
		16'h577C: out_word = 8'h57;
		16'h577D: out_word = 8'h1C;
		16'h577E: out_word = 8'hCD;
		16'h577F: out_word = 8'hFD;
		16'h5780: out_word = 8'h03;
		16'h5781: out_word = 8'h21;
		16'h5782: out_word = 8'hDD;
		16'h5783: out_word = 8'h5C;
		16'h5784: out_word = 8'h11;
		16'h5785: out_word = 8'h1A;
		16'h5786: out_word = 8'h5E;
		16'h5787: out_word = 8'h01;
		16'h5788: out_word = 8'h08;
		16'h5789: out_word = 8'h00;
		16'h578A: out_word = 8'hED;
		16'h578B: out_word = 8'hB0;
		16'h578C: out_word = 8'hCD;
		16'h578D: out_word = 8'h43;
		16'h578E: out_word = 8'h1E;
		16'h578F: out_word = 8'hC3;
		16'h5790: out_word = 8'hE1;
		16'h5791: out_word = 8'h03;
		16'h5792: out_word = 8'hFF;
		16'h5793: out_word = 8'hFF;
		16'h5794: out_word = 8'hFF;
		16'h5795: out_word = 8'hFF;
		16'h5796: out_word = 8'hFF;
		16'h5797: out_word = 8'hFF;
		16'h5798: out_word = 8'hFF;
		16'h5799: out_word = 8'hFF;
		16'h579A: out_word = 8'hFF;
		16'h579B: out_word = 8'hFF;
		16'h579C: out_word = 8'hFF;
		16'h579D: out_word = 8'hFF;
		16'h579E: out_word = 8'hFF;
		16'h579F: out_word = 8'hFF;
		16'h57A0: out_word = 8'hFF;
		16'h57A1: out_word = 8'hFF;
		16'h57A2: out_word = 8'hFF;
		16'h57A3: out_word = 8'hFF;
		16'h57A4: out_word = 8'hFF;
		16'h57A5: out_word = 8'h3A;
		16'h57A6: out_word = 8'hD3;
		16'h57A7: out_word = 8'h5C;
		16'h57A8: out_word = 8'hB7;
		16'h57A9: out_word = 8'hC8;
		16'h57AA: out_word = 8'hE5;
		16'h57AB: out_word = 8'h21;
		16'h57AC: out_word = 8'h23;
		16'h57AD: out_word = 8'h5D;
		16'h57AE: out_word = 8'h96;
		16'h57AF: out_word = 8'hE1;
		16'h57B0: out_word = 8'h30;
		16'h57B1: out_word = 8'h2B;
		16'h57B2: out_word = 8'h3A;
		16'h57B3: out_word = 8'hD3;
		16'h57B4: out_word = 8'h5C;
		16'h57B5: out_word = 8'h47;
		16'h57B6: out_word = 8'hAF;
		16'h57B7: out_word = 8'h32;
		16'h57B8: out_word = 8'hD3;
		16'h57B9: out_word = 8'h5C;
		16'h57BA: out_word = 8'hC5;
		16'h57BB: out_word = 8'h2A;
		16'h57BC: out_word = 8'hCF;
		16'h57BD: out_word = 8'h5C;
		16'h57BE: out_word = 8'hE5;
		16'h57BF: out_word = 8'hED;
		16'h57C0: out_word = 8'h5B;
		16'h57C1: out_word = 8'hD5;
		16'h57C2: out_word = 8'h5C;
		16'h57C3: out_word = 8'hCD;
		16'h57C4: out_word = 8'h3D;
		16'h57C5: out_word = 8'h1E;
		16'h57C6: out_word = 8'h2A;
		16'h57C7: out_word = 8'hF4;
		16'h57C8: out_word = 8'h5C;
		16'h57C9: out_word = 8'h22;
		16'h57CA: out_word = 8'hD5;
		16'h57CB: out_word = 8'h5C;
		16'h57CC: out_word = 8'hE1;
		16'h57CD: out_word = 8'hC1;
		16'h57CE: out_word = 8'hED;
		16'h57CF: out_word = 8'h5B;
		16'h57D0: out_word = 8'hD7;
		16'h57D1: out_word = 8'h5C;
		16'h57D2: out_word = 8'hCD;
		16'h57D3: out_word = 8'h4D;
		16'h57D4: out_word = 8'h1E;
		16'h57D5: out_word = 8'h2A;
		16'h57D6: out_word = 8'hF4;
		16'h57D7: out_word = 8'h5C;
		16'h57D8: out_word = 8'h22;
		16'h57D9: out_word = 8'hD7;
		16'h57DA: out_word = 8'h5C;
		16'h57DB: out_word = 8'h18;
		16'h57DC: out_word = 8'hC8;
		16'h57DD: out_word = 8'h32;
		16'h57DE: out_word = 8'hD3;
		16'h57DF: out_word = 8'h5C;
		16'h57E0: out_word = 8'hE5;
		16'h57E1: out_word = 8'h21;
		16'h57E2: out_word = 8'h23;
		16'h57E3: out_word = 8'h5D;
		16'h57E4: out_word = 8'h46;
		16'h57E5: out_word = 8'hE1;
		16'h57E6: out_word = 8'hAF;
		16'h57E7: out_word = 8'h18;
		16'h57E8: out_word = 8'hD1;
		16'h57E9: out_word = 8'hF5;
		16'h57EA: out_word = 8'h21;
		16'h57EB: out_word = 8'hCC;
		16'h57EC: out_word = 8'h5C;
		16'h57ED: out_word = 8'h36;
		16'h57EE: out_word = 8'h00;
		16'h57EF: out_word = 8'h79;
		16'h57F0: out_word = 8'hD6;
		16'h57F1: out_word = 8'h10;
		16'h57F2: out_word = 8'h38;
		16'h57F3: out_word = 8'h03;
		16'h57F4: out_word = 8'h34;
		16'h57F5: out_word = 8'h18;
		16'h57F6: out_word = 8'hF9;
		16'h57F7: out_word = 8'hC6;
		16'h57F8: out_word = 8'h10;
		16'h57F9: out_word = 8'h4F;
		16'h57FA: out_word = 8'hC5;
		16'h57FB: out_word = 8'hCD;
		16'h57FC: out_word = 8'hEC;
		16'h57FD: out_word = 8'h03;
		16'h57FE: out_word = 8'hC1;
		16'h57FF: out_word = 8'hF1;
		16'h5800: out_word = 8'hCD;
		16'h5801: out_word = 8'hA4;
		16'h5802: out_word = 8'h1C;
		16'h5803: out_word = 8'h11;
		16'h5804: out_word = 8'hDD;
		16'h5805: out_word = 8'h5C;
		16'h5806: out_word = 8'h01;
		16'h5807: out_word = 8'h10;
		16'h5808: out_word = 8'h00;
		16'h5809: out_word = 8'hB7;
		16'h580A: out_word = 8'h28;
		16'h580B: out_word = 8'h01;
		16'h580C: out_word = 8'hEB;
		16'h580D: out_word = 8'hED;
		16'h580E: out_word = 8'hB0;
		16'h580F: out_word = 8'hC9;
		16'h5810: out_word = 8'h3E;
		16'h5811: out_word = 8'hFF;
		16'h5812: out_word = 8'h32;
		16'h5813: out_word = 8'hF9;
		16'h5814: out_word = 8'h5C;
		16'h5815: out_word = 8'hCD;
		16'h5816: out_word = 8'h52;
		16'h5817: out_word = 8'h18;
		16'h5818: out_word = 8'hCD;
		16'h5819: out_word = 8'h36;
		16'h581A: out_word = 8'h18;
		16'h581B: out_word = 8'hCD;
		16'h581C: out_word = 8'h75;
		16'h581D: out_word = 8'h1D;
		16'h581E: out_word = 8'h3E;
		16'h581F: out_word = 8'hFF;
		16'h5820: out_word = 8'h32;
		16'h5821: out_word = 8'h10;
		16'h5822: out_word = 8'h5D;
		16'h5823: out_word = 8'h3A;
		16'h5824: out_word = 8'hF9;
		16'h5825: out_word = 8'h5C;
		16'h5826: out_word = 8'hFE;
		16'h5827: out_word = 8'hFF;
		16'h5828: out_word = 8'hCA;
		16'h5829: out_word = 8'hE1;
		16'h582A: out_word = 8'h03;
		16'h582B: out_word = 8'h3A;
		16'h582C: out_word = 8'hE5;
		16'h582D: out_word = 8'h5C;
		16'h582E: out_word = 8'hFE;
		16'h582F: out_word = 8'h42;
		16'h5830: out_word = 8'hCA;
		16'h5831: out_word = 8'h2A;
		16'h5832: out_word = 8'h01;
		16'h5833: out_word = 8'hC3;
		16'h5834: out_word = 8'hE1;
		16'h5835: out_word = 8'h03;
		16'h5836: out_word = 8'hCD;
		16'h5837: out_word = 8'h7A;
		16'h5838: out_word = 8'h18;
		16'h5839: out_word = 8'hCD;
		16'h583A: out_word = 8'h75;
		16'h583B: out_word = 8'h1D;
		16'h583C: out_word = 8'hCD;
		16'h583D: out_word = 8'hAB;
		16'h583E: out_word = 8'h18;
		16'h583F: out_word = 8'hC3;
		16'h5840: out_word = 8'h21;
		16'h5841: out_word = 8'h19;
		16'h5842: out_word = 8'h2A;
		16'h5843: out_word = 8'h5D;
		16'h5844: out_word = 8'h5C;
		16'h5845: out_word = 8'h23;
		16'h5846: out_word = 8'h7E;
		16'h5847: out_word = 8'hFE;
		16'h5848: out_word = 8'h0D;
		16'h5849: out_word = 8'hC8;
		16'h584A: out_word = 8'h3E;
		16'h584B: out_word = 8'h01;
		16'h584C: out_word = 8'h32;
		16'h584D: out_word = 8'hD6;
		16'h584E: out_word = 8'h5C;
		16'h584F: out_word = 8'hCD;
		16'h5850: out_word = 8'hEB;
		16'h5851: out_word = 8'h1D;
		16'h5852: out_word = 8'hAF;
		16'h5853: out_word = 8'h32;
		16'h5854: out_word = 8'h10;
		16'h5855: out_word = 8'h5D;
		16'h5856: out_word = 8'hC9;
		16'h5857: out_word = 8'hCD;
		16'h5858: out_word = 8'h2E;
		16'h5859: out_word = 8'h10;
		16'h585A: out_word = 8'h3E;
		16'h585B: out_word = 8'h42;
		16'h585C: out_word = 8'hB8;
		16'h585D: out_word = 8'h20;
		16'h585E: out_word = 8'h07;
		16'h585F: out_word = 8'h2A;
		16'h5860: out_word = 8'h5D;
		16'h5861: out_word = 8'h5C;
		16'h5862: out_word = 8'h2B;
		16'h5863: out_word = 8'h22;
		16'h5864: out_word = 8'h5D;
		16'h5865: out_word = 8'h5C;
		16'h5866: out_word = 8'hCD;
		16'h5867: out_word = 8'hEB;
		16'h5868: out_word = 8'h1D;
		16'h5869: out_word = 8'h2A;
		16'h586A: out_word = 8'hD9;
		16'h586B: out_word = 8'h5C;
		16'h586C: out_word = 8'h22;
		16'h586D: out_word = 8'hD7;
		16'h586E: out_word = 8'h5C;
		16'h586F: out_word = 8'h2A;
		16'h5870: out_word = 8'hDB;
		16'h5871: out_word = 8'h5C;
		16'h5872: out_word = 8'h22;
		16'h5873: out_word = 8'hD9;
		16'h5874: out_word = 8'h5C;
		16'h5875: out_word = 8'hAF;
		16'h5876: out_word = 8'h32;
		16'h5877: out_word = 8'hD6;
		16'h5878: out_word = 8'h5C;
		16'h5879: out_word = 8'hC9;
		16'h587A: out_word = 8'hCD;
		16'h587B: out_word = 8'h2B;
		16'h587C: out_word = 8'h04;
		16'h587D: out_word = 8'hCA;
		16'h587E: out_word = 8'h7B;
		16'h587F: out_word = 8'h02;
		16'h5880: out_word = 8'hCD;
		16'h5881: out_word = 8'hDF;
		16'h5882: out_word = 8'h1D;
		16'h5883: out_word = 8'hCD;
		16'h5884: out_word = 8'h72;
		16'h5885: out_word = 8'h05;
		16'h5886: out_word = 8'hC4;
		16'h5887: out_word = 8'h57;
		16'h5888: out_word = 8'h18;
		16'h5889: out_word = 8'hCD;
		16'h588A: out_word = 8'h8C;
		16'h588B: out_word = 8'h1D;
		16'h588C: out_word = 8'hFE;
		16'h588D: out_word = 8'hAF;
		16'h588E: out_word = 8'hCC;
		16'h588F: out_word = 8'h42;
		16'h5890: out_word = 8'h18;
		16'h5891: out_word = 8'hFE;
		16'h5892: out_word = 8'hE4;
		16'h5893: out_word = 8'hF5;
		16'h5894: out_word = 8'hCD;
		16'h5895: out_word = 8'h72;
		16'h5896: out_word = 8'h05;
		16'h5897: out_word = 8'hCC;
		16'h5898: out_word = 8'h2E;
		16'h5899: out_word = 8'h10;
		16'h589A: out_word = 8'hF1;
		16'h589B: out_word = 8'hCC;
		16'h589C: out_word = 8'hFC;
		16'h589D: out_word = 8'h1B;
		16'h589E: out_word = 8'hCD;
		16'h589F: out_word = 8'h75;
		16'h58A0: out_word = 8'h1D;
		16'h58A1: out_word = 8'hCD;
		16'h58A2: out_word = 8'h2F;
		16'h58A3: out_word = 8'h29;
		16'h58A4: out_word = 8'hC2;
		16'h58A5: out_word = 8'hD9;
		16'h58A6: out_word = 8'h03;
		16'h58A7: out_word = 8'hCD;
		16'h58A8: out_word = 8'h5D;
		16'h58A9: out_word = 8'h16;
		16'h58AA: out_word = 8'hC9;
		16'h58AB: out_word = 8'hCD;
		16'h58AC: out_word = 8'hCE;
		16'h58AD: out_word = 8'h33;
		16'h58AE: out_word = 8'hB7;
		16'h58AF: out_word = 8'h2A;
		16'h58B0: out_word = 8'hE6;
		16'h58B1: out_word = 8'h5C;
		16'h58B2: out_word = 8'h28;
		16'h58B3: out_word = 8'h03;
		16'h58B4: out_word = 8'h2A;
		16'h58B5: out_word = 8'hD9;
		16'h58B6: out_word = 8'h5C;
		16'h58B7: out_word = 8'hED;
		16'h58B8: out_word = 8'h5B;
		16'h58B9: out_word = 8'hEB;
		16'h58BA: out_word = 8'h5C;
		16'h58BB: out_word = 8'hFE;
		16'h58BC: out_word = 8'h03;
		16'h58BD: out_word = 8'h3A;
		16'h58BE: out_word = 8'hEA;
		16'h58BF: out_word = 8'h5C;
		16'h58C0: out_word = 8'hD5;
		16'h58C1: out_word = 8'hED;
		16'h58C2: out_word = 8'h5B;
		16'h58C3: out_word = 8'hE8;
		16'h58C4: out_word = 8'h5C;
		16'h58C5: out_word = 8'h20;
		16'h58C6: out_word = 8'h04;
		16'h58C7: out_word = 8'hED;
		16'h58C8: out_word = 8'h5B;
		16'h58C9: out_word = 8'hDB;
		16'h58CA: out_word = 8'h5C;
		16'h58CB: out_word = 8'h47;
		16'h58CC: out_word = 8'hED;
		16'h58CD: out_word = 8'h53;
		16'h58CE: out_word = 8'hDB;
		16'h58CF: out_word = 8'h5C;
		16'h58D0: out_word = 8'h3A;
		16'h58D1: out_word = 8'hE5;
		16'h58D2: out_word = 8'h5C;
		16'h58D3: out_word = 8'hFE;
		16'h58D4: out_word = 8'h43;
		16'h58D5: out_word = 8'h78;
		16'h58D6: out_word = 8'h20;
		16'h58D7: out_word = 8'h25;
		16'h58D8: out_word = 8'h78;
		16'h58D9: out_word = 8'hBA;
		16'h58DA: out_word = 8'h28;
		16'h58DB: out_word = 8'h1A;
		16'h58DC: out_word = 8'h3D;
		16'h58DD: out_word = 8'hBA;
		16'h58DE: out_word = 8'h78;
		16'h58DF: out_word = 8'h28;
		16'h58E0: out_word = 8'h15;
		16'h58E1: out_word = 8'h3A;
		16'h58E2: out_word = 8'hD6;
		16'h58E3: out_word = 8'h5C;
		16'h58E4: out_word = 8'hFE;
		16'h58E5: out_word = 8'h03;
		16'h58E6: out_word = 8'h78;
		16'h58E7: out_word = 8'h28;
		16'h58E8: out_word = 8'h0D;
		16'h58E9: out_word = 8'hAF;
		16'h58EA: out_word = 8'h32;
		16'h58EB: out_word = 8'hD6;
		16'h58EC: out_word = 8'h5C;
		16'h58ED: out_word = 8'h50;
		16'h58EE: out_word = 8'h1E;
		16'h58EF: out_word = 8'h00;
		16'h58F0: out_word = 8'hED;
		16'h58F1: out_word = 8'h53;
		16'h58F2: out_word = 8'hDB;
		16'h58F3: out_word = 8'h5C;
		16'h58F4: out_word = 8'h18;
		16'h58F5: out_word = 8'h03;
		16'h58F6: out_word = 8'hCD;
		16'h58F7: out_word = 8'h1B;
		16'h58F8: out_word = 8'h19;
		16'h58F9: out_word = 8'h78;
		16'h58FA: out_word = 8'hCD;
		16'h58FB: out_word = 8'hAC;
		16'h58FC: out_word = 8'h1E;
		16'h58FD: out_word = 8'h47;
		16'h58FE: out_word = 8'h3A;
		16'h58FF: out_word = 8'hE5;
		16'h5900: out_word = 8'h5C;
		16'h5901: out_word = 8'hFE;
		16'h5902: out_word = 8'h43;
		16'h5903: out_word = 8'hD1;
		16'h5904: out_word = 8'hC8;
		16'h5905: out_word = 8'hD5;
		16'h5906: out_word = 8'hFE;
		16'h5907: out_word = 8'h42;
		16'h5908: out_word = 8'hF5;
		16'h5909: out_word = 8'hCC;
		16'h590A: out_word = 8'h01;
		16'h590B: out_word = 8'h1A;
		16'h590C: out_word = 8'hF1;
		16'h590D: out_word = 8'hFE;
		16'h590E: out_word = 8'h44;
		16'h590F: out_word = 8'hCC;
		16'h5910: out_word = 8'h4C;
		16'h5911: out_word = 8'h1A;
		16'h5912: out_word = 8'hCD;
		16'h5913: out_word = 8'h1B;
		16'h5914: out_word = 8'h19;
		16'h5915: out_word = 8'h3A;
		16'h5916: out_word = 8'hDC;
		16'h5917: out_word = 8'h5C;
		16'h5918: out_word = 8'h47;
		16'h5919: out_word = 8'hD1;
		16'h591A: out_word = 8'hC9;
		16'h591B: out_word = 8'h3E;
		16'h591C: out_word = 8'h03;
		16'h591D: out_word = 8'h32;
		16'h591E: out_word = 8'hD6;
		16'h591F: out_word = 8'h5C;
		16'h5920: out_word = 8'hC9;
		16'h5921: out_word = 8'hCD;
		16'h5922: out_word = 8'h72;
		16'h5923: out_word = 8'h05;
		16'h5924: out_word = 8'h28;
		16'h5925: out_word = 8'h07;
		16'h5926: out_word = 8'hF5;
		16'h5927: out_word = 8'hCD;
		16'h5928: out_word = 8'h94;
		16'h5929: out_word = 8'h1A;
		16'h592A: out_word = 8'hF1;
		16'h592B: out_word = 8'hFE;
		16'h592C: out_word = 8'hFF;
		16'h592D: out_word = 8'hF5;
		16'h592E: out_word = 8'hCC;
		16'h592F: out_word = 8'h5C;
		16'h5930: out_word = 8'h19;
		16'h5931: out_word = 8'hF1;
		16'h5932: out_word = 8'h28;
		16'h5933: out_word = 8'h03;
		16'h5934: out_word = 8'hC3;
		16'h5935: out_word = 8'h4D;
		16'h5936: out_word = 8'h1E;
		16'h5937: out_word = 8'h3A;
		16'h5938: out_word = 8'hD6;
		16'h5939: out_word = 8'h5C;
		16'h593A: out_word = 8'hFE;
		16'h593B: out_word = 8'h03;
		16'h593C: out_word = 8'hCC;
		16'h593D: out_word = 8'h46;
		16'h593E: out_word = 8'h19;
		16'h593F: out_word = 8'h2A;
		16'h5940: out_word = 8'h59;
		16'h5941: out_word = 8'h5C;
		16'h5942: out_word = 8'h2B;
		16'h5943: out_word = 8'h36;
		16'h5944: out_word = 8'h80;
		16'h5945: out_word = 8'hC9;
		16'h5946: out_word = 8'h3A;
		16'h5947: out_word = 8'hF9;
		16'h5948: out_word = 8'h5C;
		16'h5949: out_word = 8'hFE;
		16'h594A: out_word = 8'hFF;
		16'h594B: out_word = 8'hC2;
		16'h594C: out_word = 8'hDE;
		16'h594D: out_word = 8'h2F;
		16'h594E: out_word = 8'h3A;
		16'h594F: out_word = 8'hDB;
		16'h5950: out_word = 8'h5C;
		16'h5951: out_word = 8'hB7;
		16'h5952: out_word = 8'hC8;
		16'h5953: out_word = 8'h4F;
		16'h5954: out_word = 8'h06;
		16'h5955: out_word = 8'h01;
		16'h5956: out_word = 8'hED;
		16'h5957: out_word = 8'h5B;
		16'h5958: out_word = 8'hF4;
		16'h5959: out_word = 8'h5C;
		16'h595A: out_word = 8'h18;
		16'h595B: out_word = 8'h0E;
		16'h595C: out_word = 8'h3A;
		16'h595D: out_word = 8'hF9;
		16'h595E: out_word = 8'h5C;
		16'h595F: out_word = 8'hFE;
		16'h5960: out_word = 8'hFF;
		16'h5961: out_word = 8'hC2;
		16'h5962: out_word = 8'h3D;
		16'h5963: out_word = 8'h1E;
		16'h5964: out_word = 8'hED;
		16'h5965: out_word = 8'h53;
		16'h5966: out_word = 8'hF4;
		16'h5967: out_word = 8'h5C;
		16'h5968: out_word = 8'h0E;
		16'h5969: out_word = 8'h00;
		16'h596A: out_word = 8'h78;
		16'h596B: out_word = 8'hB7;
		16'h596C: out_word = 8'hC8;
		16'h596D: out_word = 8'h22;
		16'h596E: out_word = 8'hD7;
		16'h596F: out_word = 8'h5C;
		16'h5970: out_word = 8'hED;
		16'h5971: out_word = 8'h53;
		16'h5972: out_word = 8'hD9;
		16'h5973: out_word = 8'h5C;
		16'h5974: out_word = 8'hC5;
		16'h5975: out_word = 8'h06;
		16'h5976: out_word = 8'h01;
		16'h5977: out_word = 8'hED;
		16'h5978: out_word = 8'h5B;
		16'h5979: out_word = 8'hD9;
		16'h597A: out_word = 8'h5C;
		16'h597B: out_word = 8'h21;
		16'h597C: out_word = 8'h25;
		16'h597D: out_word = 8'h5D;
		16'h597E: out_word = 8'hCD;
		16'h597F: out_word = 8'h3D;
		16'h5980: out_word = 8'h1E;
		16'h5981: out_word = 8'h2A;
		16'h5982: out_word = 8'hF4;
		16'h5983: out_word = 8'h5C;
		16'h5984: out_word = 8'h22;
		16'h5985: out_word = 8'hD9;
		16'h5986: out_word = 8'h5C;
		16'h5987: out_word = 8'hC1;
		16'h5988: out_word = 8'h2A;
		16'h5989: out_word = 8'hD7;
		16'h598A: out_word = 8'h5C;
		16'h598B: out_word = 8'h11;
		16'h598C: out_word = 8'h25;
		16'h598D: out_word = 8'h5D;
		16'h598E: out_word = 8'h1A;
		16'h598F: out_word = 8'hBE;
		16'h5990: out_word = 8'h20;
		16'h5991: out_word = 8'h0B;
		16'h5992: out_word = 8'h23;
		16'h5993: out_word = 8'h13;
		16'h5994: out_word = 8'h0D;
		16'h5995: out_word = 8'h20;
		16'h5996: out_word = 8'hF7;
		16'h5997: out_word = 8'h22;
		16'h5998: out_word = 8'hD7;
		16'h5999: out_word = 8'h5C;
		16'h599A: out_word = 8'h10;
		16'h599B: out_word = 8'hD8;
		16'h599C: out_word = 8'hC9;
		16'h599D: out_word = 8'h21;
		16'h599E: out_word = 8'h6B;
		16'h599F: out_word = 8'h27;
		16'h59A0: out_word = 8'h3E;
		16'h59A1: out_word = 8'h0D;
		16'h59A2: out_word = 8'hC3;
		16'h59A3: out_word = 8'h4A;
		16'h59A4: out_word = 8'h1C;
		16'h59A5: out_word = 8'h3E;
		16'h59A6: out_word = 8'hFF;
		16'h59A7: out_word = 8'h18;
		16'h59A8: out_word = 8'h02;
		16'h59A9: out_word = 8'h3E;
		16'h59AA: out_word = 8'hEE;
		16'h59AB: out_word = 8'h32;
		16'h59AC: out_word = 8'h10;
		16'h59AD: out_word = 8'h5D;
		16'h59AE: out_word = 8'hC3;
		16'h59AF: out_word = 8'h18;
		16'h59B0: out_word = 8'h18;
		16'h59B1: out_word = 8'h3E;
		16'h59B2: out_word = 8'hFF;
		16'h59B3: out_word = 8'h32;
		16'h59B4: out_word = 8'h15;
		16'h59B5: out_word = 8'h5D;
		16'h59B6: out_word = 8'hCD;
		16'h59B7: out_word = 8'h7A;
		16'h59B8: out_word = 8'h18;
		16'h59B9: out_word = 8'hCD;
		16'h59BA: out_word = 8'h75;
		16'h59BB: out_word = 8'h1D;
		16'h59BC: out_word = 8'h3A;
		16'h59BD: out_word = 8'hE5;
		16'h59BE: out_word = 8'h5C;
		16'h59BF: out_word = 8'hFE;
		16'h59C0: out_word = 8'h42;
		16'h59C1: out_word = 8'hC2;
		16'h59C2: out_word = 8'h1A;
		16'h59C3: out_word = 8'h1D;
		16'h59C4: out_word = 8'hED;
		16'h59C5: out_word = 8'h4B;
		16'h59C6: out_word = 8'hE6;
		16'h59C7: out_word = 8'h5C;
		16'h59C8: out_word = 8'hED;
		16'h59C9: out_word = 8'h43;
		16'h59CA: out_word = 8'hDB;
		16'h59CB: out_word = 8'h5C;
		16'h59CC: out_word = 8'hC5;
		16'h59CD: out_word = 8'h03;
		16'h59CE: out_word = 8'hE7;
		16'h59CF: out_word = 8'h30;
		16'h59D0: out_word = 8'h00;
		16'h59D1: out_word = 8'h36;
		16'h59D2: out_word = 8'h80;
		16'h59D3: out_word = 8'hEB;
		16'h59D4: out_word = 8'hD1;
		16'h59D5: out_word = 8'hE5;
		16'h59D6: out_word = 8'hED;
		16'h59D7: out_word = 8'h5B;
		16'h59D8: out_word = 8'hEB;
		16'h59D9: out_word = 8'h5C;
		16'h59DA: out_word = 8'hCD;
		16'h59DB: out_word = 8'h1B;
		16'h59DC: out_word = 8'h19;
		16'h59DD: out_word = 8'h3A;
		16'h59DE: out_word = 8'hDC;
		16'h59DF: out_word = 8'h5C;
		16'h59E0: out_word = 8'h47;
		16'h59E1: out_word = 8'hCD;
		16'h59E2: out_word = 8'h52;
		16'h59E3: out_word = 8'h18;
		16'h59E4: out_word = 8'hCD;
		16'h59E5: out_word = 8'h21;
		16'h59E6: out_word = 8'h19;
		16'h59E7: out_word = 8'hE1;
		16'h59E8: out_word = 8'hED;
		16'h59E9: out_word = 8'h5B;
		16'h59EA: out_word = 8'h53;
		16'h59EB: out_word = 8'h5C;
		16'h59EC: out_word = 8'hE7;
		16'h59ED: out_word = 8'hD2;
		16'h59EE: out_word = 8'h08;
		16'h59EF: out_word = 8'hC3;
		16'h59F0: out_word = 8'hE1;
		16'h59F1: out_word = 8'h03;
		16'h59F2: out_word = 8'hEB;
		16'h59F3: out_word = 8'h37;
		16'h59F4: out_word = 8'hED;
		16'h59F5: out_word = 8'h52;
		16'h59F6: out_word = 8'hD8;
		16'h59F7: out_word = 8'h11;
		16'h59F8: out_word = 8'h0A;
		16'h59F9: out_word = 8'h00;
		16'h59FA: out_word = 8'h19;
		16'h59FB: out_word = 8'h44;
		16'h59FC: out_word = 8'h4D;
		16'h59FD: out_word = 8'hE7;
		16'h59FE: out_word = 8'h05;
		16'h59FF: out_word = 8'h1F;
		16'h5A00: out_word = 8'hC9;
		16'h5A01: out_word = 8'hED;
		16'h5A02: out_word = 8'h5B;
		16'h5A03: out_word = 8'h53;
		16'h5A04: out_word = 8'h5C;
		16'h5A05: out_word = 8'h2A;
		16'h5A06: out_word = 8'h59;
		16'h5A07: out_word = 8'h5C;
		16'h5A08: out_word = 8'h2B;
		16'h5A09: out_word = 8'hE5;
		16'h5A0A: out_word = 8'hD5;
		16'h5A0B: out_word = 8'hED;
		16'h5A0C: out_word = 8'h52;
		16'h5A0D: out_word = 8'hED;
		16'h5A0E: out_word = 8'h5B;
		16'h5A0F: out_word = 8'hE6;
		16'h5A10: out_word = 8'h5C;
		16'h5A11: out_word = 8'hD5;
		16'h5A12: out_word = 8'hE5;
		16'h5A13: out_word = 8'h21;
		16'h5A14: out_word = 8'h00;
		16'h5A15: out_word = 8'h00;
		16'h5A16: out_word = 8'h3A;
		16'h5A17: out_word = 8'hF9;
		16'h5A18: out_word = 8'h5C;
		16'h5A19: out_word = 8'hFE;
		16'h5A1A: out_word = 8'hFF;
		16'h5A1B: out_word = 8'h28;
		16'h5A1C: out_word = 8'h03;
		16'h5A1D: out_word = 8'h21;
		16'h5A1E: out_word = 8'h05;
		16'h5A1F: out_word = 8'h00;
		16'h5A20: out_word = 8'h19;
		16'h5A21: out_word = 8'h22;
		16'h5A22: out_word = 8'hDB;
		16'h5A23: out_word = 8'h5C;
		16'h5A24: out_word = 8'hE1;
		16'h5A25: out_word = 8'h3A;
		16'h5A26: out_word = 8'hF9;
		16'h5A27: out_word = 8'h5C;
		16'h5A28: out_word = 8'hFE;
		16'h5A29: out_word = 8'hFF;
		16'h5A2A: out_word = 8'h20;
		16'h5A2B: out_word = 8'h05;
		16'h5A2C: out_word = 8'hD1;
		16'h5A2D: out_word = 8'hD1;
		16'h5A2E: out_word = 8'hE1;
		16'h5A2F: out_word = 8'h18;
		16'h5A30: out_word = 8'h17;
		16'h5A31: out_word = 8'hCD;
		16'h5A32: out_word = 8'hF2;
		16'h5A33: out_word = 8'h19;
		16'h5A34: out_word = 8'hC1;
		16'h5A35: out_word = 8'hD1;
		16'h5A36: out_word = 8'hE1;
		16'h5A37: out_word = 8'hC5;
		16'h5A38: out_word = 8'hE7;
		16'h5A39: out_word = 8'hE5;
		16'h5A3A: out_word = 8'h19;
		16'h5A3B: out_word = 8'hC1;
		16'h5A3C: out_word = 8'hCD;
		16'h5A3D: out_word = 8'h32;
		16'h5A3E: out_word = 8'h1E;
		16'h5A3F: out_word = 8'h23;
		16'h5A40: out_word = 8'hED;
		16'h5A41: out_word = 8'h4B;
		16'h5A42: out_word = 8'hE8;
		16'h5A43: out_word = 8'h5C;
		16'h5A44: out_word = 8'h09;
		16'h5A45: out_word = 8'h22;
		16'h5A46: out_word = 8'h4B;
		16'h5A47: out_word = 8'h5C;
		16'h5A48: out_word = 8'h2A;
		16'h5A49: out_word = 8'h53;
		16'h5A4A: out_word = 8'h5C;
		16'h5A4B: out_word = 8'hC9;
		16'h5A4C: out_word = 8'hED;
		16'h5A4D: out_word = 8'h5B;
		16'h5A4E: out_word = 8'hE8;
		16'h5A4F: out_word = 8'h5C;
		16'h5A50: out_word = 8'hED;
		16'h5A51: out_word = 8'h53;
		16'h5A52: out_word = 8'hDB;
		16'h5A53: out_word = 8'h5C;
		16'h5A54: out_word = 8'h2A;
		16'h5A55: out_word = 8'hD7;
		16'h5A56: out_word = 8'h5C;
		16'h5A57: out_word = 8'h3A;
		16'h5A58: out_word = 8'hF9;
		16'h5A59: out_word = 8'h5C;
		16'h5A5A: out_word = 8'hFE;
		16'h5A5B: out_word = 8'hFF;
		16'h5A5C: out_word = 8'hC8;
		16'h5A5D: out_word = 8'h2A;
		16'h5A5E: out_word = 8'hD9;
		16'h5A5F: out_word = 8'h5C;
		16'h5A60: out_word = 8'hE5;
		16'h5A61: out_word = 8'hCD;
		16'h5A62: out_word = 8'hF2;
		16'h5A63: out_word = 8'h19;
		16'h5A64: out_word = 8'hE1;
		16'h5A65: out_word = 8'h7C;
		16'h5A66: out_word = 8'hB5;
		16'h5A67: out_word = 8'h28;
		16'h5A68: out_word = 8'h10;
		16'h5A69: out_word = 8'h2A;
		16'h5A6A: out_word = 8'hD7;
		16'h5A6B: out_word = 8'h5C;
		16'h5A6C: out_word = 8'h2B;
		16'h5A6D: out_word = 8'h2B;
		16'h5A6E: out_word = 8'h2B;
		16'h5A6F: out_word = 8'hED;
		16'h5A70: out_word = 8'h4B;
		16'h5A71: out_word = 8'hD9;
		16'h5A72: out_word = 8'h5C;
		16'h5A73: out_word = 8'h03;
		16'h5A74: out_word = 8'h03;
		16'h5A75: out_word = 8'h03;
		16'h5A76: out_word = 8'hCD;
		16'h5A77: out_word = 8'h2E;
		16'h5A78: out_word = 8'h1E;
		16'h5A79: out_word = 8'h2A;
		16'h5A7A: out_word = 8'h59;
		16'h5A7B: out_word = 8'h5C;
		16'h5A7C: out_word = 8'h2B;
		16'h5A7D: out_word = 8'hED;
		16'h5A7E: out_word = 8'h4B;
		16'h5A7F: out_word = 8'hE8;
		16'h5A80: out_word = 8'h5C;
		16'h5A81: out_word = 8'hC5;
		16'h5A82: out_word = 8'h03;
		16'h5A83: out_word = 8'h03;
		16'h5A84: out_word = 8'h03;
		16'h5A85: out_word = 8'hCD;
		16'h5A86: out_word = 8'h32;
		16'h5A87: out_word = 8'h1E;
		16'h5A88: out_word = 8'h23;
		16'h5A89: out_word = 8'h3A;
		16'h5A8A: out_word = 8'hD2;
		16'h5A8B: out_word = 8'h5C;
		16'h5A8C: out_word = 8'h77;
		16'h5A8D: out_word = 8'h23;
		16'h5A8E: out_word = 8'hD1;
		16'h5A8F: out_word = 8'h73;
		16'h5A90: out_word = 8'h23;
		16'h5A91: out_word = 8'h72;
		16'h5A92: out_word = 8'h23;
		16'h5A93: out_word = 8'hC9;
		16'h5A94: out_word = 8'h3A;
		16'h5A95: out_word = 8'hD9;
		16'h5A96: out_word = 8'h5C;
		16'h5A97: out_word = 8'h48;
		16'h5A98: out_word = 8'h47;
		16'h5A99: out_word = 8'h79;
		16'h5A9A: out_word = 8'hB8;
		16'h5A9B: out_word = 8'h38;
		16'h5A9C: out_word = 8'h19;
		16'h5A9D: out_word = 8'h78;
		16'h5A9E: out_word = 8'hB7;
		16'h5A9F: out_word = 8'hCA;
		16'h5AA0: out_word = 8'h1A;
		16'h5AA1: out_word = 8'h1D;
		16'h5AA2: out_word = 8'h05;
		16'h5AA3: out_word = 8'h28;
		16'h5AA4: out_word = 8'h0B;
		16'h5AA5: out_word = 8'h3E;
		16'h5AA6: out_word = 8'h10;
		16'h5AA7: out_word = 8'h1C;
		16'h5AA8: out_word = 8'hBB;
		16'h5AA9: out_word = 8'h20;
		16'h5AAA: out_word = 8'h03;
		16'h5AAB: out_word = 8'h1E;
		16'h5AAC: out_word = 8'h00;
		16'h5AAD: out_word = 8'h14;
		16'h5AAE: out_word = 8'h10;
		16'h5AAF: out_word = 8'hF7;
		16'h5AB0: out_word = 8'h06;
		16'h5AB1: out_word = 8'h01;
		16'h5AB2: out_word = 8'h2A;
		16'h5AB3: out_word = 8'hD7;
		16'h5AB4: out_word = 8'h5C;
		16'h5AB5: out_word = 8'hC9;
		16'h5AB6: out_word = 8'h21;
		16'h5AB7: out_word = 8'hED;
		16'h5AB8: out_word = 8'h29;
		16'h5AB9: out_word = 8'h3E;
		16'h5ABA: out_word = 8'h05;
		16'h5ABB: out_word = 8'hC3;
		16'h5ABC: out_word = 8'h4A;
		16'h5ABD: out_word = 8'h1C;
		16'h5ABE: out_word = 8'hCD;
		16'h5ABF: out_word = 8'h2F;
		16'h5AC0: out_word = 8'h29;
		16'h5AC1: out_word = 8'hCC;
		16'h5AC2: out_word = 8'h43;
		16'h5AC3: out_word = 8'h33;
		16'h5AC4: out_word = 8'hCD;
		16'h5AC5: out_word = 8'hFD;
		16'h5AC6: out_word = 8'h03;
		16'h5AC7: out_word = 8'h3A;
		16'h5AC8: out_word = 8'h09;
		16'h5AC9: out_word = 8'h5E;
		16'h5ACA: out_word = 8'hFE;
		16'h5ACB: out_word = 8'h80;
		16'h5ACC: out_word = 8'hCA;
		16'h5ACD: out_word = 8'h23;
		16'h5ACE: out_word = 8'h27;
		16'h5ACF: out_word = 8'hC9;
		16'h5AD0: out_word = 8'hCD;
		16'h5AD1: out_word = 8'h52;
		16'h5AD2: out_word = 8'h18;
		16'h5AD3: out_word = 8'h21;
		16'h5AD4: out_word = 8'h00;
		16'h5AD5: out_word = 8'h00;
		16'h5AD6: out_word = 8'h22;
		16'h5AD7: out_word = 8'hD1;
		16'h5AD8: out_word = 8'h5C;
		16'h5AD9: out_word = 8'hCD;
		16'h5ADA: out_word = 8'hDF;
		16'h5ADB: out_word = 8'h1D;
		16'h5ADC: out_word = 8'hCD;
		16'h5ADD: out_word = 8'h8C;
		16'h5ADE: out_word = 8'h1D;
		16'h5ADF: out_word = 8'hFE;
		16'h5AE0: out_word = 8'hAF;
		16'h5AE1: out_word = 8'h28;
		16'h5AE2: out_word = 8'h56;
		16'h5AE3: out_word = 8'hFE;
		16'h5AE4: out_word = 8'hCA;
		16'h5AE5: out_word = 8'h20;
		16'h5AE6: out_word = 8'h11;
		16'h5AE7: out_word = 8'hCD;
		16'h5AE8: out_word = 8'h0B;
		16'h5AE9: out_word = 8'h1E;
		16'h5AEA: out_word = 8'hCD;
		16'h5AEB: out_word = 8'h75;
		16'h5AEC: out_word = 8'h1D;
		16'h5AED: out_word = 8'h2A;
		16'h5AEE: out_word = 8'hDB;
		16'h5AEF: out_word = 8'h5C;
		16'h5AF0: out_word = 8'h22;
		16'h5AF1: out_word = 8'hD1;
		16'h5AF2: out_word = 8'h5C;
		16'h5AF3: out_word = 8'h21;
		16'h5AF4: out_word = 8'hE5;
		16'h5AF5: out_word = 8'h5C;
		16'h5AF6: out_word = 8'h18;
		16'h5AF7: out_word = 8'h27;
		16'h5AF8: out_word = 8'hFE;
		16'h5AF9: out_word = 8'hAA;
		16'h5AFA: out_word = 8'h20;
		16'h5AFB: out_word = 8'h11;
		16'h5AFC: out_word = 8'h21;
		16'h5AFD: out_word = 8'h00;
		16'h5AFE: out_word = 8'h40;
		16'h5AFF: out_word = 8'h22;
		16'h5B00: out_word = 8'hD7;
		16'h5B01: out_word = 8'h5C;
		16'h5B02: out_word = 8'h21;
		16'h5B03: out_word = 8'h00;
		16'h5B04: out_word = 8'h1B;
		16'h5B05: out_word = 8'h22;
		16'h5B06: out_word = 8'hD9;
		16'h5B07: out_word = 8'h5C;
		16'h5B08: out_word = 8'h22;
		16'h5B09: out_word = 8'hDB;
		16'h5B0A: out_word = 8'h5C;
		16'h5B0B: out_word = 8'h18;
		16'h5B0C: out_word = 8'h3B;
		16'h5B0D: out_word = 8'hCD;
		16'h5B0E: out_word = 8'h75;
		16'h5B0F: out_word = 8'h1D;
		16'h5B10: out_word = 8'hCD;
		16'h5B11: out_word = 8'h8C;
		16'h5B12: out_word = 8'h1D;
		16'h5B13: out_word = 8'h21;
		16'h5B14: out_word = 8'hE5;
		16'h5B15: out_word = 8'h5C;
		16'h5B16: out_word = 8'hFE;
		16'h5B17: out_word = 8'hE4;
		16'h5B18: out_word = 8'h28;
		16'h5B19: out_word = 8'h12;
		16'h5B1A: out_word = 8'hFE;
		16'h5B1B: out_word = 8'h0D;
		16'h5B1C: out_word = 8'hC2;
		16'h5B1D: out_word = 8'h1A;
		16'h5B1E: out_word = 8'h1D;
		16'h5B1F: out_word = 8'h36;
		16'h5B20: out_word = 8'h42;
		16'h5B21: out_word = 8'hCD;
		16'h5B22: out_word = 8'hBE;
		16'h5B23: out_word = 8'h1A;
		16'h5B24: out_word = 8'hCD;
		16'h5B25: out_word = 8'h1C;
		16'h5B26: out_word = 8'h1E;
		16'h5B27: out_word = 8'hCD;
		16'h5B28: out_word = 8'hDE;
		16'h5B29: out_word = 8'h1B;
		16'h5B2A: out_word = 8'h18;
		16'h5B2B: out_word = 8'h27;
		16'h5B2C: out_word = 8'h36;
		16'h5B2D: out_word = 8'h44;
		16'h5B2E: out_word = 8'hCD;
		16'h5B2F: out_word = 8'hBE;
		16'h5B30: out_word = 8'h1A;
		16'h5B31: out_word = 8'hCD;
		16'h5B32: out_word = 8'h0F;
		16'h5B33: out_word = 8'h1C;
		16'h5B34: out_word = 8'h30;
		16'h5B35: out_word = 8'h1D;
		16'h5B36: out_word = 8'hDA;
		16'h5B37: out_word = 8'h1A;
		16'h5B38: out_word = 8'h1D;
		16'h5B39: out_word = 8'hCD;
		16'h5B3A: out_word = 8'hE5;
		16'h5B3B: out_word = 8'h1D;
		16'h5B3C: out_word = 8'h2A;
		16'h5B3D: out_word = 8'hD9;
		16'h5B3E: out_word = 8'h5C;
		16'h5B3F: out_word = 8'h22;
		16'h5B40: out_word = 8'hD7;
		16'h5B41: out_word = 8'h5C;
		16'h5B42: out_word = 8'h2A;
		16'h5B43: out_word = 8'hDB;
		16'h5B44: out_word = 8'h5C;
		16'h5B45: out_word = 8'h22;
		16'h5B46: out_word = 8'hD9;
		16'h5B47: out_word = 8'h5C;
		16'h5B48: out_word = 8'hCD;
		16'h5B49: out_word = 8'h75;
		16'h5B4A: out_word = 8'h1D;
		16'h5B4B: out_word = 8'h3E;
		16'h5B4C: out_word = 8'h43;
		16'h5B4D: out_word = 8'h32;
		16'h5B4E: out_word = 8'hE5;
		16'h5B4F: out_word = 8'h5C;
		16'h5B50: out_word = 8'hCD;
		16'h5B51: out_word = 8'hBE;
		16'h5B52: out_word = 8'h1A;
		16'h5B53: out_word = 8'hCD;
		16'h5B54: out_word = 8'hF5;
		16'h5B55: out_word = 8'h33;
		16'h5B56: out_word = 8'hC3;
		16'h5B57: out_word = 8'h69;
		16'h5B58: out_word = 8'h05;
		16'h5B59: out_word = 8'h2A;
		16'h5B5A: out_word = 8'hD7;
		16'h5B5B: out_word = 8'h5C;
		16'h5B5C: out_word = 8'h22;
		16'h5B5D: out_word = 8'hE6;
		16'h5B5E: out_word = 8'h5C;
		16'h5B5F: out_word = 8'hEB;
		16'h5B60: out_word = 8'h2A;
		16'h5B61: out_word = 8'hD9;
		16'h5B62: out_word = 8'h5C;
		16'h5B63: out_word = 8'h7D;
		16'h5B64: out_word = 8'hB4;
		16'h5B65: out_word = 8'hCA;
		16'h5B66: out_word = 8'h1A;
		16'h5B67: out_word = 8'h1D;
		16'h5B68: out_word = 8'h7D;
		16'h5B69: out_word = 8'hB7;
		16'h5B6A: out_word = 8'h28;
		16'h5B6B: out_word = 8'h01;
		16'h5B6C: out_word = 8'h24;
		16'h5B6D: out_word = 8'h7C;
		16'h5B6E: out_word = 8'h32;
		16'h5B6F: out_word = 8'hEA;
		16'h5B70: out_word = 8'h5C;
		16'h5B71: out_word = 8'h5F;
		16'h5B72: out_word = 8'h16;
		16'h5B73: out_word = 8'h00;
		16'h5B74: out_word = 8'h2A;
		16'h5B75: out_word = 8'h0A;
		16'h5B76: out_word = 8'h5E;
		16'h5B77: out_word = 8'hED;
		16'h5B78: out_word = 8'h52;
		16'h5B79: out_word = 8'hDA;
		16'h5B7A: out_word = 8'h45;
		16'h5B7B: out_word = 8'h1C;
		16'h5B7C: out_word = 8'hE5;
		16'h5B7D: out_word = 8'h2A;
		16'h5B7E: out_word = 8'h59;
		16'h5B7F: out_word = 8'h5C;
		16'h5B80: out_word = 8'h36;
		16'h5B81: out_word = 8'hAA;
		16'h5B82: out_word = 8'h23;
		16'h5B83: out_word = 8'hED;
		16'h5B84: out_word = 8'h5B;
		16'h5B85: out_word = 8'hD1;
		16'h5B86: out_word = 8'h5C;
		16'h5B87: out_word = 8'h73;
		16'h5B88: out_word = 8'h23;
		16'h5B89: out_word = 8'h72;
		16'h5B8A: out_word = 8'h2A;
		16'h5B8B: out_word = 8'hDB;
		16'h5B8C: out_word = 8'h5C;
		16'h5B8D: out_word = 8'h22;
		16'h5B8E: out_word = 8'hE8;
		16'h5B8F: out_word = 8'h5C;
		16'h5B90: out_word = 8'h2A;
		16'h5B91: out_word = 8'h06;
		16'h5B92: out_word = 8'h5E;
		16'h5B93: out_word = 8'h22;
		16'h5B94: out_word = 8'hEB;
		16'h5B95: out_word = 8'h5C;
		16'h5B96: out_word = 8'hEB;
		16'h5B97: out_word = 8'h2A;
		16'h5B98: out_word = 8'hE6;
		16'h5B99: out_word = 8'h5C;
		16'h5B9A: out_word = 8'h3A;
		16'h5B9B: out_word = 8'hEA;
		16'h5B9C: out_word = 8'h5C;
		16'h5B9D: out_word = 8'h47;
		16'h5B9E: out_word = 8'hCD;
		16'h5B9F: out_word = 8'h4D;
		16'h5BA0: out_word = 8'h1E;
		16'h5BA1: out_word = 8'h2A;
		16'h5BA2: out_word = 8'hF4;
		16'h5BA3: out_word = 8'h5C;
		16'h5BA4: out_word = 8'hE5;
		16'h5BA5: out_word = 8'hCD;
		16'h5BA6: out_word = 8'hFD;
		16'h5BA7: out_word = 8'h03;
		16'h5BA8: out_word = 8'hE1;
		16'h5BA9: out_word = 8'h22;
		16'h5BAA: out_word = 8'h06;
		16'h5BAB: out_word = 8'h5E;
		16'h5BAC: out_word = 8'hE1;
		16'h5BAD: out_word = 8'h22;
		16'h5BAE: out_word = 8'h0A;
		16'h5BAF: out_word = 8'h5E;
		16'h5BB0: out_word = 8'h21;
		16'h5BB1: out_word = 8'h09;
		16'h5BB2: out_word = 8'h5E;
		16'h5BB3: out_word = 8'h7E;
		16'h5BB4: out_word = 8'h32;
		16'h5BB5: out_word = 8'h1E;
		16'h5BB6: out_word = 8'h5D;
		16'h5BB7: out_word = 8'h34;
		16'h5BB8: out_word = 8'hE5;
		16'h5BB9: out_word = 8'hCD;
		16'h5BBA: out_word = 8'h43;
		16'h5BBB: out_word = 8'h1E;
		16'h5BBC: out_word = 8'hE1;
		16'h5BBD: out_word = 8'h4E;
		16'h5BBE: out_word = 8'h0D;
		16'h5BBF: out_word = 8'h3A;
		16'h5BC0: out_word = 8'hE5;
		16'h5BC1: out_word = 8'h5C;
		16'h5BC2: out_word = 8'hFE;
		16'h5BC3: out_word = 8'h42;
		16'h5BC4: out_word = 8'hCC;
		16'h5BC5: out_word = 8'hC8;
		16'h5BC6: out_word = 8'h1B;
		16'h5BC7: out_word = 8'hC9;
		16'h5BC8: out_word = 8'h2A;
		16'h5BC9: out_word = 8'h59;
		16'h5BCA: out_word = 8'h5C;
		16'h5BCB: out_word = 8'hED;
		16'h5BCC: out_word = 8'h5B;
		16'h5BCD: out_word = 8'h53;
		16'h5BCE: out_word = 8'h5C;
		16'h5BCF: out_word = 8'h37;
		16'h5BD0: out_word = 8'hED;
		16'h5BD1: out_word = 8'h52;
		16'h5BD2: out_word = 8'h22;
		16'h5BD3: out_word = 8'hE6;
		16'h5BD4: out_word = 8'h5C;
		16'h5BD5: out_word = 8'h2A;
		16'h5BD6: out_word = 8'h4B;
		16'h5BD7: out_word = 8'h5C;
		16'h5BD8: out_word = 8'hED;
		16'h5BD9: out_word = 8'h52;
		16'h5BDA: out_word = 8'h22;
		16'h5BDB: out_word = 8'hE8;
		16'h5BDC: out_word = 8'h5C;
		16'h5BDD: out_word = 8'hC9;
		16'h5BDE: out_word = 8'h2A;
		16'h5BDF: out_word = 8'h4B;
		16'h5BE0: out_word = 8'h5C;
		16'h5BE1: out_word = 8'hED;
		16'h5BE2: out_word = 8'h5B;
		16'h5BE3: out_word = 8'h53;
		16'h5BE4: out_word = 8'h5C;
		16'h5BE5: out_word = 8'hED;
		16'h5BE6: out_word = 8'h52;
		16'h5BE7: out_word = 8'h22;
		16'h5BE8: out_word = 8'hDB;
		16'h5BE9: out_word = 8'h5C;
		16'h5BEA: out_word = 8'h2A;
		16'h5BEB: out_word = 8'h53;
		16'h5BEC: out_word = 8'h5C;
		16'h5BED: out_word = 8'h22;
		16'h5BEE: out_word = 8'hD7;
		16'h5BEF: out_word = 8'h5C;
		16'h5BF0: out_word = 8'h2A;
		16'h5BF1: out_word = 8'h59;
		16'h5BF2: out_word = 8'h5C;
		16'h5BF3: out_word = 8'h23;
		16'h5BF4: out_word = 8'h23;
		16'h5BF5: out_word = 8'h23;
		16'h5BF6: out_word = 8'hED;
		16'h5BF7: out_word = 8'h52;
		16'h5BF8: out_word = 8'h22;
		16'h5BF9: out_word = 8'hD9;
		16'h5BFA: out_word = 8'h5C;
		16'h5BFB: out_word = 8'hC9;
		16'h5BFC: out_word = 8'hCD;
		16'h5BFD: out_word = 8'h1B;
		16'h5BFE: out_word = 8'h1C;
		16'h5BFF: out_word = 8'hD0;
		16'h5C00: out_word = 8'h21;
		16'h5C01: out_word = 8'h00;
		16'h5C02: out_word = 8'h00;
		16'h5C03: out_word = 8'h22;
		16'h5C04: out_word = 8'hD9;
		16'h5C05: out_word = 8'h5C;
		16'h5C06: out_word = 8'h3A;
		16'h5C07: out_word = 8'hF9;
		16'h5C08: out_word = 8'h5C;
		16'h5C09: out_word = 8'hFE;
		16'h5C0A: out_word = 8'hFF;
		16'h5C0B: out_word = 8'hC0;
		16'h5C0C: out_word = 8'hC3;
		16'h5C0D: out_word = 8'h13;
		16'h5C0E: out_word = 8'h1C;
		16'h5C0F: out_word = 8'hCD;
		16'h5C10: out_word = 8'h1B;
		16'h5C11: out_word = 8'h1C;
		16'h5C12: out_word = 8'hD0;
		16'h5C13: out_word = 8'h3E;
		16'h5C14: out_word = 8'h0E;
		16'h5C15: out_word = 8'h21;
		16'h5C16: out_word = 8'hDD;
		16'h5C17: out_word = 8'h27;
		16'h5C18: out_word = 8'hC3;
		16'h5C19: out_word = 8'h4A;
		16'h5C1A: out_word = 8'h1C;
		16'h5C1B: out_word = 8'hCD;
		16'h5C1C: out_word = 8'h2A;
		16'h5C1D: out_word = 8'h1E;
		16'h5C1E: out_word = 8'hCD;
		16'h5C1F: out_word = 8'h9B;
		16'h5C20: out_word = 8'h1D;
		16'h5C21: out_word = 8'hCB;
		16'h5C22: out_word = 8'hF9;
		16'h5C23: out_word = 8'h79;
		16'h5C24: out_word = 8'h32;
		16'h5C25: out_word = 8'hD2;
		16'h5C26: out_word = 8'h5C;
		16'h5C27: out_word = 8'h30;
		16'h5C28: out_word = 8'h02;
		16'h5C29: out_word = 8'h37;
		16'h5C2A: out_word = 8'hC9;
		16'h5C2B: out_word = 8'h20;
		16'h5C2C: out_word = 8'hFC;
		16'h5C2D: out_word = 8'h23;
		16'h5C2E: out_word = 8'h5E;
		16'h5C2F: out_word = 8'h23;
		16'h5C30: out_word = 8'h56;
		16'h5C31: out_word = 8'h23;
		16'h5C32: out_word = 8'h22;
		16'h5C33: out_word = 8'hD7;
		16'h5C34: out_word = 8'h5C;
		16'h5C35: out_word = 8'hED;
		16'h5C36: out_word = 8'h53;
		16'h5C37: out_word = 8'hDB;
		16'h5C38: out_word = 8'h5C;
		16'h5C39: out_word = 8'hED;
		16'h5C3A: out_word = 8'h53;
		16'h5C3B: out_word = 8'hD9;
		16'h5C3C: out_word = 8'h5C;
		16'h5C3D: out_word = 8'hCD;
		16'h5C3E: out_word = 8'h2A;
		16'h5C3F: out_word = 8'h1E;
		16'h5C40: out_word = 8'hFE;
		16'h5C41: out_word = 8'h29;
		16'h5C42: out_word = 8'h20;
		16'h5C43: out_word = 8'hE7;
		16'h5C44: out_word = 8'hC9;
		16'h5C45: out_word = 8'h21;
		16'h5C46: out_word = 8'hBB;
		16'h5C47: out_word = 8'h29;
		16'h5C48: out_word = 8'h3E;
		16'h5C49: out_word = 8'h03;
		16'h5C4A: out_word = 8'hCD;
		16'h5C4B: out_word = 8'hC3;
		16'h5C4C: out_word = 8'h03;
		16'h5C4D: out_word = 8'hC3;
		16'h5C4E: out_word = 8'hD3;
		16'h5C4F: out_word = 8'h01;
		16'h5C50: out_word = 8'h21;
		16'h5C51: out_word = 8'hC5;
		16'h5C52: out_word = 8'h29;
		16'h5C53: out_word = 8'h3E;
		16'h5C54: out_word = 8'h02;
		16'h5C55: out_word = 8'h18;
		16'h5C56: out_word = 8'hF3;
		16'h5C57: out_word = 8'h21;
		16'h5C58: out_word = 8'hDD;
		16'h5C59: out_word = 8'h5C;
		16'h5C5A: out_word = 8'h06;
		16'h5C5B: out_word = 8'h08;
		16'h5C5C: out_word = 8'h36;
		16'h5C5D: out_word = 8'h20;
		16'h5C5E: out_word = 8'h23;
		16'h5C5F: out_word = 8'h10;
		16'h5C60: out_word = 8'hFB;
		16'h5C61: out_word = 8'hCD;
		16'h5C62: out_word = 8'h31;
		16'h5C63: out_word = 8'h05;
		16'h5C64: out_word = 8'hEB;
		16'h5C65: out_word = 8'hCD;
		16'h5C66: out_word = 8'h81;
		16'h5C67: out_word = 8'h1C;
		16'h5C68: out_word = 8'h79;
		16'h5C69: out_word = 8'hB0;
		16'h5C6A: out_word = 8'hCA;
		16'h5C6B: out_word = 8'h1A;
		16'h5C6C: out_word = 8'h1D;
		16'h5C6D: out_word = 8'hFE;
		16'h5C6E: out_word = 8'h09;
		16'h5C6F: out_word = 8'h38;
		16'h5C70: out_word = 8'h02;
		16'h5C71: out_word = 8'h0E;
		16'h5C72: out_word = 8'h08;
		16'h5C73: out_word = 8'h7E;
		16'h5C74: out_word = 8'hFE;
		16'h5C75: out_word = 8'h20;
		16'h5C76: out_word = 8'hDA;
		16'h5C77: out_word = 8'h1A;
		16'h5C78: out_word = 8'h1D;
		16'h5C79: out_word = 8'h11;
		16'h5C7A: out_word = 8'hDD;
		16'h5C7B: out_word = 8'h5C;
		16'h5C7C: out_word = 8'hC5;
		16'h5C7D: out_word = 8'hED;
		16'h5C7E: out_word = 8'hB0;
		16'h5C7F: out_word = 8'hC1;
		16'h5C80: out_word = 8'hC9;
		16'h5C81: out_word = 8'h23;
		16'h5C82: out_word = 8'h7E;
		16'h5C83: out_word = 8'hFE;
		16'h5C84: out_word = 8'h3A;
		16'h5C85: out_word = 8'h20;
		16'h5C86: out_word = 8'h11;
		16'h5C87: out_word = 8'h2B;
		16'h5C88: out_word = 8'h7E;
		16'h5C89: out_word = 8'hCD;
		16'h5C8A: out_word = 8'h24;
		16'h5C8B: out_word = 8'h05;
		16'h5C8C: out_word = 8'hC5;
		16'h5C8D: out_word = 8'hE5;
		16'h5C8E: out_word = 8'hCD;
		16'h5C8F: out_word = 8'hCB;
		16'h5C90: out_word = 8'h3D;
		16'h5C91: out_word = 8'hE1;
		16'h5C92: out_word = 8'hC1;
		16'h5C93: out_word = 8'h0B;
		16'h5C94: out_word = 8'h0B;
		16'h5C95: out_word = 8'h23;
		16'h5C96: out_word = 8'h23;
		16'h5C97: out_word = 8'hC9;
		16'h5C98: out_word = 8'h2B;
		16'h5C99: out_word = 8'h3A;
		16'h5C9A: out_word = 8'h19;
		16'h5C9B: out_word = 8'h5D;
		16'h5C9C: out_word = 8'hC5;
		16'h5C9D: out_word = 8'hE5;
		16'h5C9E: out_word = 8'hCD;
		16'h5C9F: out_word = 8'hCB;
		16'h5CA0: out_word = 8'h3D;
		16'h5CA1: out_word = 8'hE1;
		16'h5CA2: out_word = 8'hC1;
		16'h5CA3: out_word = 8'hC9;
		16'h5CA4: out_word = 8'h69;
		16'h5CA5: out_word = 8'h26;
		16'h5CA6: out_word = 8'h00;
		16'h5CA7: out_word = 8'h29;
		16'h5CA8: out_word = 8'h29;
		16'h5CA9: out_word = 8'h29;
		16'h5CAA: out_word = 8'h29;
		16'h5CAB: out_word = 8'h01;
		16'h5CAC: out_word = 8'h25;
		16'h5CAD: out_word = 8'h5D;
		16'h5CAE: out_word = 8'h09;
		16'h5CAF: out_word = 8'hC9;
		16'h5CB0: out_word = 8'hCD;
		16'h5CB1: out_word = 8'h57;
		16'h5CB2: out_word = 8'h1C;
		16'h5CB3: out_word = 8'hCD;
		16'h5CB4: out_word = 8'hE8;
		16'h5CB5: out_word = 8'h03;
		16'h5CB6: out_word = 8'h06;
		16'h5CB7: out_word = 8'h80;
		16'h5CB8: out_word = 8'h0E;
		16'h5CB9: out_word = 8'h00;
		16'h5CBA: out_word = 8'hC5;
		16'h5CBB: out_word = 8'hCD;
		16'h5CBC: out_word = 8'hA4;
		16'h5CBD: out_word = 8'h1C;
		16'h5CBE: out_word = 8'hCD;
		16'h5CBF: out_word = 8'h0C;
		16'h5CC0: out_word = 8'h05;
		16'h5CC1: out_word = 8'hC1;
		16'h5CC2: out_word = 8'hC5;
		16'h5CC3: out_word = 8'h79;
		16'h5CC4: out_word = 8'hFE;
		16'h5CC5: out_word = 8'h10;
		16'h5CC6: out_word = 8'h20;
		16'h5CC7: out_word = 8'h05;
		16'h5CC8: out_word = 8'hC1;
		16'h5CC9: out_word = 8'h0E;
		16'h5CCA: out_word = 8'h00;
		16'h5CCB: out_word = 8'h18;
		16'h5CCC: out_word = 8'hED;
		16'h5CCD: out_word = 8'h11;
		16'h5CCE: out_word = 8'hDD;
		16'h5CCF: out_word = 8'h5C;
		16'h5CD0: out_word = 8'h3A;
		16'h5CD1: out_word = 8'h06;
		16'h5CD2: out_word = 8'h5D;
		16'h5CD3: out_word = 8'h47;
		16'h5CD4: out_word = 8'hAF;
		16'h5CD5: out_word = 8'hBE;
		16'h5CD6: out_word = 8'h20;
		16'h5CD7: out_word = 8'h03;
		16'h5CD8: out_word = 8'hC1;
		16'h5CD9: out_word = 8'h18;
		16'h5CDA: out_word = 8'h09;
		16'h5CDB: out_word = 8'hCD;
		16'h5CDC: out_word = 8'h13;
		16'h5CDD: out_word = 8'h27;
		16'h5CDE: out_word = 8'hC1;
		16'h5CDF: out_word = 8'h28;
		16'h5CE0: out_word = 8'h06;
		16'h5CE1: out_word = 8'h0C;
		16'h5CE2: out_word = 8'h10;
		16'h5CE3: out_word = 8'hD6;
		16'h5CE4: out_word = 8'hF6;
		16'h5CE5: out_word = 8'hFF;
		16'h5CE6: out_word = 8'hC9;
		16'h5CE7: out_word = 8'h3E;
		16'h5CE8: out_word = 8'h80;
		16'h5CE9: out_word = 8'h90;
		16'h5CEA: out_word = 8'h4F;
		16'h5CEB: out_word = 8'h32;
		16'h5CEC: out_word = 8'h1E;
		16'h5CED: out_word = 8'h5D;
		16'h5CEE: out_word = 8'hAF;
		16'h5CEF: out_word = 8'hC8;
		16'h5CF0: out_word = 8'hCD;
		16'h5CF1: out_word = 8'hB3;
		16'h5CF2: out_word = 8'h1C;
		16'h5CF3: out_word = 8'h21;
		16'h5CF4: out_word = 8'h0F;
		16'h5CF5: out_word = 8'h5D;
		16'h5CF6: out_word = 8'h71;
		16'h5CF7: out_word = 8'hC8;
		16'h5CF8: out_word = 8'h36;
		16'h5CF9: out_word = 8'hFF;
		16'h5CFA: out_word = 8'hC9;
		16'h5CFB: out_word = 8'hCD;
		16'h5CFC: out_word = 8'h75;
		16'h5CFD: out_word = 8'h1D;
		16'h5CFE: out_word = 8'hCD;
		16'h5CFF: out_word = 8'hE5;
		16'h5D00: out_word = 8'h20;
		16'h5D01: out_word = 8'hFD;
		16'h5D02: out_word = 8'hCB;
		16'h5D03: out_word = 8'h01;
		16'h5D04: out_word = 8'h9E;
		16'h5D05: out_word = 8'hCD;
		16'h5D06: out_word = 8'h32;
		16'h5D07: out_word = 8'h02;
		16'h5D08: out_word = 8'hED;
		16'h5D09: out_word = 8'h7B;
		16'h5D0A: out_word = 8'h1C;
		16'h5D0B: out_word = 8'h5D;
		16'h5D0C: out_word = 8'hD9;
		16'h5D0D: out_word = 8'h21;
		16'h5D0E: out_word = 8'h58;
		16'h5D0F: out_word = 8'h27;
		16'h5D10: out_word = 8'hD9;
		16'h5D11: out_word = 8'h2B;
		16'h5D12: out_word = 8'h3E;
		16'h5D13: out_word = 8'h12;
		16'h5D14: out_word = 8'hBE;
		16'h5D15: out_word = 8'hC0;
		16'h5D16: out_word = 8'h2B;
		16'h5D17: out_word = 8'hC3;
		16'h5D18: out_word = 8'h35;
		16'h5D19: out_word = 8'h02;
		16'h5D1A: out_word = 8'hFD;
		16'h5D1B: out_word = 8'hCB;
		16'h5D1C: out_word = 8'h00;
		16'h5D1D: out_word = 8'h7E;
		16'h5D1E: out_word = 8'h28;
		16'h5D1F: out_word = 8'h05;
		16'h5D20: out_word = 8'h3E;
		16'h5D21: out_word = 8'h0B;
		16'h5D22: out_word = 8'h32;
		16'h5D23: out_word = 8'h3A;
		16'h5D24: out_word = 8'h5C;
		16'h5D25: out_word = 8'h3C;
		16'h5D26: out_word = 8'h21;
		16'h5D27: out_word = 8'hB2;
		16'h5D28: out_word = 8'h29;
		16'h5D29: out_word = 8'hCD;
		16'h5D2A: out_word = 8'hC3;
		16'h5D2B: out_word = 8'h03;
		16'h5D2C: out_word = 8'hC3;
		16'h5D2D: out_word = 8'hD3;
		16'h5D2E: out_word = 8'h01;
		16'h5D2F: out_word = 8'h3A;
		16'h5D30: out_word = 8'h3A;
		16'h5D31: out_word = 8'h5C;
		16'h5D32: out_word = 8'h21;
		16'h5D33: out_word = 8'hCA;
		16'h5D34: out_word = 8'h27;
		16'h5D35: out_word = 8'hFE;
		16'h5D36: out_word = 8'h14;
		16'h5D37: out_word = 8'h28;
		16'h5D38: out_word = 8'hF0;
		16'h5D39: out_word = 8'hFE;
		16'h5D3A: out_word = 8'h0C;
		16'h5D3B: out_word = 8'h28;
		16'h5D3C: out_word = 8'hEC;
		16'h5D3D: out_word = 8'h21;
		16'h5D3E: out_word = 8'hD2;
		16'h5D3F: out_word = 8'h27;
		16'h5D40: out_word = 8'hFE;
		16'h5D41: out_word = 8'h03;
		16'h5D42: out_word = 8'h28;
		16'h5D43: out_word = 8'hE5;
		16'h5D44: out_word = 8'h21;
		16'h5D45: out_word = 8'hDD;
		16'h5D46: out_word = 8'h27;
		16'h5D47: out_word = 8'hFE;
		16'h5D48: out_word = 8'h01;
		16'h5D49: out_word = 8'h28;
		16'h5D4A: out_word = 8'hDE;
		16'h5D4B: out_word = 8'h18;
		16'h5D4C: out_word = 8'hCD;
		16'h5D4D: out_word = 8'hCD;
		16'h5D4E: out_word = 8'h52;
		16'h5D4F: out_word = 8'h18;
		16'h5D50: out_word = 8'hCD;
		16'h5D51: out_word = 8'h36;
		16'h5D52: out_word = 8'h18;
		16'h5D53: out_word = 8'hCD;
		16'h5D54: out_word = 8'h75;
		16'h5D55: out_word = 8'h1D;
		16'h5D56: out_word = 8'h2A;
		16'h5D57: out_word = 8'hE6;
		16'h5D58: out_word = 8'h5C;
		16'h5D59: out_word = 8'h3A;
		16'h5D5A: out_word = 8'hE5;
		16'h5D5B: out_word = 8'h5C;
		16'h5D5C: out_word = 8'hFE;
		16'h5D5D: out_word = 8'h42;
		16'h5D5E: out_word = 8'hCA;
		16'h5D5F: out_word = 8'h2A;
		16'h5D60: out_word = 8'h01;
		16'h5D61: out_word = 8'hE5;
		16'h5D62: out_word = 8'hC9;
		16'h5D63: out_word = 8'h21;
		16'h5D64: out_word = 8'h0E;
		16'h5D65: out_word = 8'h5D;
		16'h5D66: out_word = 8'h7E;
		16'h5D67: out_word = 8'hFE;
		16'h5D68: out_word = 8'hFF;
		16'h5D69: out_word = 8'h36;
		16'h5D6A: out_word = 8'h00;
		16'h5D6B: out_word = 8'hC0;
		16'h5D6C: out_word = 8'hE7;
		16'h5D6D: out_word = 8'hBF;
		16'h5D6E: out_word = 8'h16;
		16'h5D6F: out_word = 8'hC9;
		16'h5D70: out_word = 8'hFD;
		16'h5D71: out_word = 8'hCB;
		16'h5D72: out_word = 8'h01;
		16'h5D73: out_word = 8'h7E;
		16'h5D74: out_word = 8'hC9;
		16'h5D75: out_word = 8'hCD;
		16'h5D76: out_word = 8'h70;
		16'h5D77: out_word = 8'h1D;
		16'h5D78: out_word = 8'hC0;
		16'h5D79: out_word = 8'hE1;
		16'h5D7A: out_word = 8'hC9;
		16'h5D7B: out_word = 8'hCD;
		16'h5D7C: out_word = 8'h2A;
		16'h5D7D: out_word = 8'h1E;
		16'h5D7E: out_word = 8'hCD;
		16'h5D7F: out_word = 8'hC1;
		16'h5D80: out_word = 8'h1D;
		16'h5D81: out_word = 8'h18;
		16'h5D82: out_word = 8'hED;
		16'h5D83: out_word = 8'hAF;
		16'h5D84: out_word = 8'hE7;
		16'h5D85: out_word = 8'h01;
		16'h5D86: out_word = 8'h16;
		16'h5D87: out_word = 8'hC9;
		16'h5D88: out_word = 8'h3E;
		16'h5D89: out_word = 8'h02;
		16'h5D8A: out_word = 8'h18;
		16'h5D8B: out_word = 8'hF8;
		16'h5D8C: out_word = 8'hE7;
		16'h5D8D: out_word = 8'h18;
		16'h5D8E: out_word = 8'h00;
		16'h5D8F: out_word = 8'hC9;
		16'h5D90: out_word = 8'hCD;
		16'h5D91: out_word = 8'h83;
		16'h5D92: out_word = 8'h1D;
		16'h5D93: out_word = 8'hE7;
		16'h5D94: out_word = 8'h2C;
		16'h5D95: out_word = 8'h0F;
		16'h5D96: out_word = 8'hC9;
		16'h5D97: out_word = 8'hE7;
		16'h5D98: out_word = 8'h6B;
		16'h5D99: out_word = 8'h0D;
		16'h5D9A: out_word = 8'hC9;
		16'h5D9B: out_word = 8'hE7;
		16'h5D9C: out_word = 8'hB2;
		16'h5D9D: out_word = 8'h28;
		16'h5D9E: out_word = 8'hC9;
		16'h5D9F: out_word = 8'hE7;
		16'h5DA0: out_word = 8'h6E;
		16'h5DA1: out_word = 8'h0D;
		16'h5DA2: out_word = 8'hC9;
		16'h5DA3: out_word = 8'h4F;
		16'h5DA4: out_word = 8'h06;
		16'h5DA5: out_word = 8'h00;
		16'h5DA6: out_word = 8'hC3;
		16'h5DA7: out_word = 8'hA9;
		16'h5DA8: out_word = 8'h1D;
		16'h5DA9: out_word = 8'hC5;
		16'h5DAA: out_word = 8'hCD;
		16'h5DAB: out_word = 8'hF1;
		16'h5DAC: out_word = 8'h20;
		16'h5DAD: out_word = 8'hC1;
		16'h5DAE: out_word = 8'hE7;
		16'h5DAF: out_word = 8'h1B;
		16'h5DB0: out_word = 8'h1A;
		16'h5DB1: out_word = 8'hCD;
		16'h5DB2: out_word = 8'hF1;
		16'h5DB3: out_word = 8'h20;
		16'h5DB4: out_word = 8'hC9;
		16'h5DB5: out_word = 8'hE7;
		16'h5DB6: out_word = 8'hF1;
		16'h5DB7: out_word = 8'h2B;
		16'h5DB8: out_word = 8'hC9;
		16'h5DB9: out_word = 8'hE7;
		16'h5DBA: out_word = 8'h99;
		16'h5DBB: out_word = 8'h1E;
		16'h5DBC: out_word = 8'hC9;
		16'h5DBD: out_word = 8'hE7;
		16'h5DBE: out_word = 8'h8C;
		16'h5DBF: out_word = 8'h1C;
		16'h5DC0: out_word = 8'hC9;
		16'h5DC1: out_word = 8'hE7;
		16'h5DC2: out_word = 8'h82;
		16'h5DC3: out_word = 8'h1C;
		16'h5DC4: out_word = 8'hC9;
		16'h5DC5: out_word = 8'h2A;
		16'h5DC6: out_word = 8'h11;
		16'h5DC7: out_word = 8'h5D;
		16'h5DC8: out_word = 8'h23;
		16'h5DC9: out_word = 8'h22;
		16'h5DCA: out_word = 8'h5D;
		16'h5DCB: out_word = 8'h5C;
		16'h5DCC: out_word = 8'hC9;
		16'h5DCD: out_word = 8'hCD;
		16'h5DCE: out_word = 8'hDF;
		16'h5DCF: out_word = 8'h1D;
		16'h5DD0: out_word = 8'hCD;
		16'h5DD1: out_word = 8'h8C;
		16'h5DD2: out_word = 8'h1D;
		16'h5DD3: out_word = 8'hFE;
		16'h5DD4: out_word = 8'h2C;
		16'h5DD5: out_word = 8'hC2;
		16'h5DD6: out_word = 8'h1A;
		16'h5DD7: out_word = 8'h1D;
		16'h5DD8: out_word = 8'hCD;
		16'h5DD9: out_word = 8'h2A;
		16'h5DDA: out_word = 8'h1E;
		16'h5DDB: out_word = 8'hCD;
		16'h5DDC: out_word = 8'hBD;
		16'h5DDD: out_word = 8'h1D;
		16'h5DDE: out_word = 8'hC9;
		16'h5DDF: out_word = 8'hCD;
		16'h5DE0: out_word = 8'hC5;
		16'h5DE1: out_word = 8'h1D;
		16'h5DE2: out_word = 8'hC3;
		16'h5DE3: out_word = 8'hBD;
		16'h5DE4: out_word = 8'h1D;
		16'h5DE5: out_word = 8'hCD;
		16'h5DE6: out_word = 8'h8C;
		16'h5DE7: out_word = 8'h1D;
		16'h5DE8: out_word = 8'hFE;
		16'h5DE9: out_word = 8'hAF;
		16'h5DEA: out_word = 8'hC0;
		16'h5DEB: out_word = 8'hCD;
		16'h5DEC: out_word = 8'h7B;
		16'h5DED: out_word = 8'h1D;
		16'h5DEE: out_word = 8'h28;
		16'h5DEF: out_word = 8'h0B;
		16'h5DF0: out_word = 8'hCD;
		16'h5DF1: out_word = 8'hB9;
		16'h5DF2: out_word = 8'h1D;
		16'h5DF3: out_word = 8'hED;
		16'h5DF4: out_word = 8'h43;
		16'h5DF5: out_word = 8'hD9;
		16'h5DF6: out_word = 8'h5C;
		16'h5DF7: out_word = 8'hED;
		16'h5DF8: out_word = 8'h43;
		16'h5DF9: out_word = 8'hDB;
		16'h5DFA: out_word = 8'h5C;
		16'h5DFB: out_word = 8'hCD;
		16'h5DFC: out_word = 8'h8C;
		16'h5DFD: out_word = 8'h1D;
		16'h5DFE: out_word = 8'hFE;
		16'h5DFF: out_word = 8'h2C;
		16'h5E00: out_word = 8'h28;
		16'h5E01: out_word = 8'h09;
		16'h5E02: out_word = 8'hFE;
		16'h5E03: out_word = 8'h0D;
		16'h5E04: out_word = 8'hC2;
		16'h5E05: out_word = 8'h1A;
		16'h5E06: out_word = 8'h1D;
		16'h5E07: out_word = 8'hCD;
		16'h5E08: out_word = 8'h75;
		16'h5E09: out_word = 8'h1D;
		16'h5E0A: out_word = 8'hC9;
		16'h5E0B: out_word = 8'hCD;
		16'h5E0C: out_word = 8'h7B;
		16'h5E0D: out_word = 8'h1D;
		16'h5E0E: out_word = 8'hC8;
		16'h5E0F: out_word = 8'hCD;
		16'h5E10: out_word = 8'hB9;
		16'h5E11: out_word = 8'h1D;
		16'h5E12: out_word = 8'hED;
		16'h5E13: out_word = 8'h43;
		16'h5E14: out_word = 8'hDB;
		16'h5E15: out_word = 8'h5C;
		16'h5E16: out_word = 8'h3E;
		16'h5E17: out_word = 8'h03;
		16'h5E18: out_word = 8'h32;
		16'h5E19: out_word = 8'hD6;
		16'h5E1A: out_word = 8'h5C;
		16'h5E1B: out_word = 8'hC9;
		16'h5E1C: out_word = 8'h2A;
		16'h5E1D: out_word = 8'h11;
		16'h5E1E: out_word = 8'h5D;
		16'h5E1F: out_word = 8'hE7;
		16'h5E20: out_word = 8'hA7;
		16'h5E21: out_word = 8'h11;
		16'h5E22: out_word = 8'hC9;
		16'h5E23: out_word = 8'h2A;
		16'h5E24: out_word = 8'h61;
		16'h5E25: out_word = 8'h5C;
		16'h5E26: out_word = 8'hE7;
		16'h5E27: out_word = 8'h30;
		16'h5E28: out_word = 8'h00;
		16'h5E29: out_word = 8'hC9;
		16'h5E2A: out_word = 8'hE7;
		16'h5E2B: out_word = 8'h20;
		16'h5E2C: out_word = 8'h00;
		16'h5E2D: out_word = 8'hC9;
		16'h5E2E: out_word = 8'hE7;
		16'h5E2F: out_word = 8'hE8;
		16'h5E30: out_word = 8'h19;
		16'h5E31: out_word = 8'hC9;
		16'h5E32: out_word = 8'hE7;
		16'h5E33: out_word = 8'h55;
		16'h5E34: out_word = 8'h16;
		16'h5E35: out_word = 8'hC9;
		16'h5E36: out_word = 8'hCD;
		16'h5E37: out_word = 8'hB2;
		16'h5E38: out_word = 8'h3E;
		16'h5E39: out_word = 8'h7C;
		16'h5E3A: out_word = 8'hD3;
		16'h5E3B: out_word = 8'h3F;
		16'h5E3C: out_word = 8'hC9;
		16'h5E3D: out_word = 8'hAF;
		16'h5E3E: out_word = 8'h18;
		16'h5E3F: out_word = 8'h24;
		16'h5E40: out_word = 8'hCD;
		16'h5E41: out_word = 8'h6B;
		16'h5E42: out_word = 8'h16;
		16'h5E43: out_word = 8'hED;
		16'h5E44: out_word = 8'h5B;
		16'h5E45: out_word = 8'hF4;
		16'h5E46: out_word = 8'h5C;
		16'h5E47: out_word = 8'h1B;
		16'h5E48: out_word = 8'h06;
		16'h5E49: out_word = 8'h01;
		16'h5E4A: out_word = 8'h21;
		16'h5E4B: out_word = 8'h25;
		16'h5E4C: out_word = 8'h5D;
		16'h5E4D: out_word = 8'hE5;
		16'h5E4E: out_word = 8'hD5;
		16'h5E4F: out_word = 8'hCD;
		16'h5E50: out_word = 8'h11;
		16'h5E51: out_word = 8'h3E;
		16'h5E52: out_word = 8'hCB;
		16'h5E53: out_word = 8'h7E;
		16'h5E54: out_word = 8'h28;
		16'h5E55: out_word = 8'h0A;
		16'h5E56: out_word = 8'hCB;
		16'h5E57: out_word = 8'h46;
		16'h5E58: out_word = 8'h20;
		16'h5E59: out_word = 8'h06;
		16'h5E5A: out_word = 8'h21;
		16'h5E5B: out_word = 8'hD8;
		16'h5E5C: out_word = 8'h29;
		16'h5E5D: out_word = 8'hC3;
		16'h5E5E: out_word = 8'h29;
		16'h5E5F: out_word = 8'h1D;
		16'h5E60: out_word = 8'hD1;
		16'h5E61: out_word = 8'hE1;
		16'h5E62: out_word = 8'h3E;
		16'h5E63: out_word = 8'hFF;
		16'h5E64: out_word = 8'h32;
		16'h5E65: out_word = 8'hCE;
		16'h5E66: out_word = 8'h5C;
		16'h5E67: out_word = 8'hED;
		16'h5E68: out_word = 8'h53;
		16'h5E69: out_word = 8'hF4;
		16'h5E6A: out_word = 8'h5C;
		16'h5E6B: out_word = 8'hC5;
		16'h5E6C: out_word = 8'hE5;
		16'h5E6D: out_word = 8'hC3;
		16'h5E6E: out_word = 8'h00;
		16'h5E6F: out_word = 8'h38;
		16'h5E70: out_word = 8'hE1;
		16'h5E71: out_word = 8'hC1;
		16'h5E72: out_word = 8'hAF;
		16'h5E73: out_word = 8'hB0;
		16'h5E74: out_word = 8'hC8;
		16'h5E75: out_word = 8'hC5;
		16'h5E76: out_word = 8'hE5;
		16'h5E77: out_word = 8'hCD;
		16'h5E78: out_word = 8'h06;
		16'h5E79: out_word = 8'h3F;
		16'h5E7A: out_word = 8'h3A;
		16'h5E7B: out_word = 8'hF4;
		16'h5E7C: out_word = 8'h5C;
		16'h5E7D: out_word = 8'hCD;
		16'h5E7E: out_word = 8'h02;
		16'h5E7F: out_word = 8'h3F;
		16'h5E80: out_word = 8'h3A;
		16'h5E81: out_word = 8'hF5;
		16'h5E82: out_word = 8'h5C;
		16'h5E83: out_word = 8'hCD;
		16'h5E84: out_word = 8'h63;
		16'h5E85: out_word = 8'h3E;
		16'h5E86: out_word = 8'h3A;
		16'h5E87: out_word = 8'hCE;
		16'h5E88: out_word = 8'h5C;
		16'h5E89: out_word = 8'hB7;
		16'h5E8A: out_word = 8'hF5;
		16'h5E8B: out_word = 8'hCC;
		16'h5E8C: out_word = 8'h0E;
		16'h5E8D: out_word = 8'h3F;
		16'h5E8E: out_word = 8'hF1;
		16'h5E8F: out_word = 8'hC4;
		16'h5E90: out_word = 8'h0A;
		16'h5E91: out_word = 8'h3F;
		16'h5E92: out_word = 8'hE1;
		16'h5E93: out_word = 8'h11;
		16'h5E94: out_word = 8'h00;
		16'h5E95: out_word = 8'h01;
		16'h5E96: out_word = 8'h19;
		16'h5E97: out_word = 8'hE5;
		16'h5E98: out_word = 8'h3E;
		16'h5E99: out_word = 8'h10;
		16'h5E9A: out_word = 8'h21;
		16'h5E9B: out_word = 8'hF4;
		16'h5E9C: out_word = 8'h5C;
		16'h5E9D: out_word = 8'h34;
		16'h5E9E: out_word = 8'hBE;
		16'h5E9F: out_word = 8'h20;
		16'h5EA0: out_word = 8'h06;
		16'h5EA1: out_word = 8'h36;
		16'h5EA2: out_word = 8'h00;
		16'h5EA3: out_word = 8'h21;
		16'h5EA4: out_word = 8'hF5;
		16'h5EA5: out_word = 8'h5C;
		16'h5EA6: out_word = 8'h34;
		16'h5EA7: out_word = 8'hE1;
		16'h5EA8: out_word = 8'hC1;
		16'h5EA9: out_word = 8'h10;
		16'h5EAA: out_word = 8'hCA;
		16'h5EAB: out_word = 8'hC9;
		16'h5EAC: out_word = 8'hE5;
		16'h5EAD: out_word = 8'h67;
		16'h5EAE: out_word = 8'h2E;
		16'h5EAF: out_word = 8'h00;
		16'h5EB0: out_word = 8'hE5;
		16'h5EB1: out_word = 8'hED;
		16'h5EB2: out_word = 8'h52;
		16'h5EB3: out_word = 8'hDC;
		16'h5EB4: out_word = 8'hBC;
		16'h5EB5: out_word = 8'h1E;
		16'h5EB6: out_word = 8'hE1;
		16'h5EB7: out_word = 8'h7C;
		16'h5EB8: out_word = 8'hE1;
		16'h5EB9: out_word = 8'hD8;
		16'h5EBA: out_word = 8'h7A;
		16'h5EBB: out_word = 8'hC9;
		16'h5EBC: out_word = 8'hAF;
		16'h5EBD: out_word = 8'h32;
		16'h5EBE: out_word = 8'hD6;
		16'h5EBF: out_word = 8'h5C;
		16'h5EC0: out_word = 8'h37;
		16'h5EC1: out_word = 8'hC9;
		16'h5EC2: out_word = 8'h21;
		16'h5EC3: out_word = 8'hFF;
		16'h5EC4: out_word = 8'hFF;
		16'h5EC5: out_word = 8'h22;
		16'h5EC6: out_word = 8'hD7;
		16'h5EC7: out_word = 8'h5C;
		16'h5EC8: out_word = 8'h22;
		16'h5EC9: out_word = 8'hD9;
		16'h5ECA: out_word = 8'h5C;
		16'h5ECB: out_word = 8'h22;
		16'h5ECC: out_word = 8'hD1;
		16'h5ECD: out_word = 8'h5C;
		16'h5ECE: out_word = 8'hCD;
		16'h5ECF: out_word = 8'h2B;
		16'h5ED0: out_word = 8'h04;
		16'h5ED1: out_word = 8'hCA;
		16'h5ED2: out_word = 8'h1A;
		16'h5ED3: out_word = 8'h1D;
		16'h5ED4: out_word = 8'hCD;
		16'h5ED5: out_word = 8'hDF;
		16'h5ED6: out_word = 8'h1D;
		16'h5ED7: out_word = 8'hCD;
		16'h5ED8: out_word = 8'h75;
		16'h5ED9: out_word = 8'h1D;
		16'h5EDA: out_word = 8'hCD;
		16'h5EDB: out_word = 8'h21;
		16'h5EDC: out_word = 8'h39;
		16'h5EDD: out_word = 8'hCD;
		16'h5EDE: out_word = 8'h78;
		16'h5EDF: out_word = 8'h33;
		16'h5EE0: out_word = 8'hE6;
		16'h5EE1: out_word = 8'h80;
		16'h5EE2: out_word = 8'h3E;
		16'h5EE3: out_word = 8'h28;
		16'h5EE4: out_word = 8'h28;
		16'h5EE5: out_word = 8'h02;
		16'h5EE6: out_word = 8'h3E;
		16'h5EE7: out_word = 8'h50;
		16'h5EE8: out_word = 8'h32;
		16'h5EE9: out_word = 8'hD7;
		16'h5EEA: out_word = 8'h5C;
		16'h5EEB: out_word = 8'hCD;
		16'h5EEC: out_word = 8'h98;
		16'h5EED: out_word = 8'h3D;
		16'h5EEE: out_word = 8'hCD;
		16'h5EEF: out_word = 8'hF6;
		16'h5EF0: out_word = 8'h1F;
		16'h5EF1: out_word = 8'hCD;
		16'h5EF2: out_word = 8'hA0;
		16'h5EF3: out_word = 8'h3E;
		16'h5EF4: out_word = 8'hCD;
		16'h5EF5: out_word = 8'hBC;
		16'h5EF6: out_word = 8'h1E;
		16'h5EF7: out_word = 8'h3A;
		16'h5EF8: out_word = 8'hDD;
		16'h5EF9: out_word = 8'h5C;
		16'h5EFA: out_word = 8'hFE;
		16'h5EFB: out_word = 8'h24;
		16'h5EFC: out_word = 8'h28;
		16'h5EFD: out_word = 8'h1D;
		16'h5EFE: out_word = 8'h18;
		16'h5EFF: out_word = 8'h16;
		16'h5F00: out_word = 8'hFF;
		16'h5F01: out_word = 8'hFF;
		16'h5F02: out_word = 8'hFF;
		16'h5F03: out_word = 8'hFF;
		16'h5F04: out_word = 8'hFF;
		16'h5F05: out_word = 8'hFF;
		16'h5F06: out_word = 8'hFF;
		16'h5F07: out_word = 8'hFF;
		16'h5F08: out_word = 8'hFF;
		16'h5F09: out_word = 8'hFF;
		16'h5F0A: out_word = 8'hFF;
		16'h5F0B: out_word = 8'hFF;
		16'h5F0C: out_word = 8'hFF;
		16'h5F0D: out_word = 8'hFF;
		16'h5F0E: out_word = 8'hFF;
		16'h5F0F: out_word = 8'hFF;
		16'h5F10: out_word = 8'hFF;
		16'h5F11: out_word = 8'hFF;
		16'h5F12: out_word = 8'hFF;
		16'h5F13: out_word = 8'hFF;
		16'h5F14: out_word = 8'hFF;
		16'h5F15: out_word = 8'hFF;
		16'h5F16: out_word = 8'h3E;
		16'h5F17: out_word = 8'h80;
		16'h5F18: out_word = 8'h32;
		16'h5F19: out_word = 8'hDA;
		16'h5F1A: out_word = 8'h5C;
		16'h5F1B: out_word = 8'hCD;
		16'h5F1C: out_word = 8'h4C;
		16'h5F1D: out_word = 8'h33;
		16'h5F1E: out_word = 8'h21;
		16'h5F1F: out_word = 8'h25;
		16'h5F20: out_word = 8'h5D;
		16'h5F21: out_word = 8'h36;
		16'h5F22: out_word = 8'h00;
		16'h5F23: out_word = 8'h11;
		16'h5F24: out_word = 8'h26;
		16'h5F25: out_word = 8'h5D;
		16'h5F26: out_word = 8'h01;
		16'h5F27: out_word = 8'hFF;
		16'h5F28: out_word = 8'h00;
		16'h5F29: out_word = 8'hED;
		16'h5F2A: out_word = 8'hB0;
		16'h5F2B: out_word = 8'h01;
		16'h5F2C: out_word = 8'hD7;
		16'h5F2D: out_word = 8'h5C;
		16'h5F2E: out_word = 8'h11;
		16'h5F2F: out_word = 8'hDA;
		16'h5F30: out_word = 8'h5C;
		16'h5F31: out_word = 8'h0A;
		16'h5F32: out_word = 8'hFE;
		16'h5F33: out_word = 8'h50;
		16'h5F34: out_word = 8'h28;
		16'h5F35: out_word = 8'h13;
		16'h5F36: out_word = 8'h1A;
		16'h5F37: out_word = 8'hFE;
		16'h5F38: out_word = 8'h80;
		16'h5F39: out_word = 8'h28;
		16'h5F3A: out_word = 8'h07;
		16'h5F3B: out_word = 8'h3E;
		16'h5F3C: out_word = 8'h19;
		16'h5F3D: out_word = 8'h21;
		16'h5F3E: out_word = 8'h70;
		16'h5F3F: out_word = 8'h02;
		16'h5F40: out_word = 8'h18;
		16'h5F41: out_word = 8'h13;
		16'h5F42: out_word = 8'h3E;
		16'h5F43: out_word = 8'h17;
		16'h5F44: out_word = 8'h21;
		16'h5F45: out_word = 8'hF0;
		16'h5F46: out_word = 8'h04;
		16'h5F47: out_word = 8'h18;
		16'h5F48: out_word = 8'h0C;
		16'h5F49: out_word = 8'h1A;
		16'h5F4A: out_word = 8'hFE;
		16'h5F4B: out_word = 8'h80;
		16'h5F4C: out_word = 8'h3E;
		16'h5F4D: out_word = 8'h18;
		16'h5F4E: out_word = 8'h20;
		16'h5F4F: out_word = 8'hF4;
		16'h5F50: out_word = 8'h3E;
		16'h5F51: out_word = 8'h16;
		16'h5F52: out_word = 8'h21;
		16'h5F53: out_word = 8'hF0;
		16'h5F54: out_word = 8'h09;
		16'h5F55: out_word = 8'h32;
		16'h5F56: out_word = 8'h08;
		16'h5F57: out_word = 8'h5E;
		16'h5F58: out_word = 8'h22;
		16'h5F59: out_word = 8'h0A;
		16'h5F5A: out_word = 8'h5E;
		16'h5F5B: out_word = 8'h3E;
		16'h5F5C: out_word = 8'h01;
		16'h5F5D: out_word = 8'h32;
		16'h5F5E: out_word = 8'h07;
		16'h5F5F: out_word = 8'h5E;
		16'h5F60: out_word = 8'h3E;
		16'h5F61: out_word = 8'h10;
		16'h5F62: out_word = 8'h32;
		16'h5F63: out_word = 8'h0C;
		16'h5F64: out_word = 8'h5E;
		16'h5F65: out_word = 8'h21;
		16'h5F66: out_word = 8'h0F;
		16'h5F67: out_word = 8'h5E;
		16'h5F68: out_word = 8'h11;
		16'h5F69: out_word = 8'h10;
		16'h5F6A: out_word = 8'h5E;
		16'h5F6B: out_word = 8'h01;
		16'h5F6C: out_word = 8'h08;
		16'h5F6D: out_word = 8'h00;
		16'h5F6E: out_word = 8'h36;
		16'h5F6F: out_word = 8'h20;
		16'h5F70: out_word = 8'hED;
		16'h5F71: out_word = 8'hB0;
		16'h5F72: out_word = 8'h21;
		16'h5F73: out_word = 8'hDD;
		16'h5F74: out_word = 8'h5C;
		16'h5F75: out_word = 8'h11;
		16'h5F76: out_word = 8'h1A;
		16'h5F77: out_word = 8'h5E;
		16'h5F78: out_word = 8'h01;
		16'h5F79: out_word = 8'h08;
		16'h5F7A: out_word = 8'h00;
		16'h5F7B: out_word = 8'hED;
		16'h5F7C: out_word = 8'hB0;
		16'h5F7D: out_word = 8'hCD;
		16'h5F7E: out_word = 8'hEB;
		16'h5F7F: out_word = 8'h1F;
		16'h5F80: out_word = 8'h06;
		16'h5F81: out_word = 8'h01;
		16'h5F82: out_word = 8'h11;
		16'h5F83: out_word = 8'h08;
		16'h5F84: out_word = 8'h00;
		16'h5F85: out_word = 8'h21;
		16'h5F86: out_word = 8'h25;
		16'h5F87: out_word = 8'h5D;
		16'h5F88: out_word = 8'hCD;
		16'h5F89: out_word = 8'h62;
		16'h5F8A: out_word = 8'h1E;
		16'h5F8B: out_word = 8'h3A;
		16'h5F8C: out_word = 8'hD6;
		16'h5F8D: out_word = 8'h5C;
		16'h5F8E: out_word = 8'hF5;
		16'h5F8F: out_word = 8'hAF;
		16'h5F90: out_word = 8'h32;
		16'h5F91: out_word = 8'hE5;
		16'h5F92: out_word = 8'h5C;
		16'h5F93: out_word = 8'h2A;
		16'h5F94: out_word = 8'h0A;
		16'h5F95: out_word = 8'h5E;
		16'h5F96: out_word = 8'h22;
		16'h5F97: out_word = 8'hD7;
		16'h5F98: out_word = 8'h5C;
		16'h5F99: out_word = 8'h21;
		16'h5F9A: out_word = 8'hDD;
		16'h5F9B: out_word = 8'h5C;
		16'h5F9C: out_word = 8'hDF;
		16'h5F9D: out_word = 8'h3E;
		16'h5F9E: out_word = 8'h0D;
		16'h5F9F: out_word = 8'hD7;
		16'h5FA0: out_word = 8'h2A;
		16'h5FA1: out_word = 8'hD7;
		16'h5FA2: out_word = 8'h5C;
		16'h5FA3: out_word = 8'hF1;
		16'h5FA4: out_word = 8'hE5;
		16'h5FA5: out_word = 8'h16;
		16'h5FA6: out_word = 8'h00;
		16'h5FA7: out_word = 8'h5F;
		16'h5FA8: out_word = 8'hED;
		16'h5FA9: out_word = 8'h52;
		16'h5FAA: out_word = 8'h44;
		16'h5FAB: out_word = 8'h4D;
		16'h5FAC: out_word = 8'hCD;
		16'h5FAD: out_word = 8'hA9;
		16'h5FAE: out_word = 8'h1D;
		16'h5FAF: out_word = 8'h3E;
		16'h5FB0: out_word = 8'h2F;
		16'h5FB1: out_word = 8'hD7;
		16'h5FB2: out_word = 8'hC1;
		16'h5FB3: out_word = 8'hCD;
		16'h5FB4: out_word = 8'hA9;
		16'h5FB5: out_word = 8'h1D;
		16'h5FB6: out_word = 8'hC3;
		16'h5FB7: out_word = 8'h33;
		16'h5FB8: out_word = 8'h08;
		16'h5FB9: out_word = 8'h01;
		16'h5FBA: out_word = 8'h09;
		16'h5FBB: out_word = 8'h02;
		16'h5FBC: out_word = 8'h0A;
		16'h5FBD: out_word = 8'h03;
		16'h5FBE: out_word = 8'h0B;
		16'h5FBF: out_word = 8'h04;
		16'h5FC0: out_word = 8'h0C;
		16'h5FC1: out_word = 8'h05;
		16'h5FC2: out_word = 8'h0D;
		16'h5FC3: out_word = 8'h06;
		16'h5FC4: out_word = 8'h0E;
		16'h5FC5: out_word = 8'h07;
		16'h5FC6: out_word = 8'h0F;
		16'h5FC7: out_word = 8'h08;
		16'h5FC8: out_word = 8'h10;
		16'h5FC9: out_word = 8'h01;
		16'h5FCA: out_word = 8'hCD;
		16'h5FCB: out_word = 8'h08;
		16'h5FCC: out_word = 8'h3E;
		16'h5FCD: out_word = 8'hF6;
		16'h5FCE: out_word = 8'h11;
		16'h5FCF: out_word = 8'h47;
		16'h5FD0: out_word = 8'h3E;
		16'h5FD1: out_word = 8'h32;
		16'h5FD2: out_word = 8'hCD;
		16'h5FD3: out_word = 8'h44;
		16'h5FD4: out_word = 8'h3E;
		16'h5FD5: out_word = 8'h3E;
		16'h5FD6: out_word = 8'h02;
		16'h5FD7: out_word = 8'hCD;
		16'h5FD8: out_word = 8'h44;
		16'h5FD9: out_word = 8'h3E;
		16'h5FDA: out_word = 8'hCD;
		16'h5FDB: out_word = 8'hFD;
		16'h5FDC: out_word = 8'h3D;
		16'h5FDD: out_word = 8'hDB;
		16'h5FDE: out_word = 8'h1F;
		16'h5FDF: out_word = 8'hE6;
		16'h5FE0: out_word = 8'h04;
		16'h5FE1: out_word = 8'h3E;
		16'h5FE2: out_word = 8'h50;
		16'h5FE3: out_word = 8'h28;
		16'h5FE4: out_word = 8'h02;
		16'h5FE5: out_word = 8'h3E;
		16'h5FE6: out_word = 8'h28;
		16'h5FE7: out_word = 8'h32;
		16'h5FE8: out_word = 8'hD7;
		16'h5FE9: out_word = 8'h5C;
		16'h5FEA: out_word = 8'hC9;
		16'h5FEB: out_word = 8'h3A;
		16'h5FEC: out_word = 8'h16;
		16'h5FED: out_word = 8'h5D;
		16'h5FEE: out_word = 8'hF6;
		16'h5FEF: out_word = 8'h3C;
		16'h5FF0: out_word = 8'h32;
		16'h5FF1: out_word = 8'h16;
		16'h5FF2: out_word = 8'h5D;
		16'h5FF3: out_word = 8'hD3;
		16'h5FF4: out_word = 8'hFF;
		16'h5FF5: out_word = 8'hC9;
		16'h5FF6: out_word = 8'h3A;
		16'h5FF7: out_word = 8'h16;
		16'h5FF8: out_word = 8'h5D;
		16'h5FF9: out_word = 8'hE6;
		16'h5FFA: out_word = 8'h6F;
		16'h5FFB: out_word = 8'h18;
		16'h5FFC: out_word = 8'hF3;
		16'h5FFD: out_word = 8'hF3;
		16'h5FFE: out_word = 8'h3E;
		16'h5FFF: out_word = 8'hF4;
		16'h6000: out_word = 8'hD3;
		16'h6001: out_word = 8'h1F;
		16'h6002: out_word = 8'h2A;
		16'h6003: out_word = 8'hE6;
		16'h6004: out_word = 8'h5C;
		16'h6005: out_word = 8'h0E;
		16'h6006: out_word = 8'h7F;
		16'h6007: out_word = 8'h06;
		16'h6008: out_word = 8'h0A;
		16'h6009: out_word = 8'h16;
		16'h600A: out_word = 8'h4E;
		16'h600B: out_word = 8'hCD;
		16'h600C: out_word = 8'hB1;
		16'h600D: out_word = 8'h20;
		16'h600E: out_word = 8'h06;
		16'h600F: out_word = 8'h0C;
		16'h6010: out_word = 8'h16;
		16'h6011: out_word = 8'h00;
		16'h6012: out_word = 8'hCD;
		16'h6013: out_word = 8'hB1;
		16'h6014: out_word = 8'h20;
		16'h6015: out_word = 8'h06;
		16'h6016: out_word = 8'h03;
		16'h6017: out_word = 8'h16;
		16'h6018: out_word = 8'hF5;
		16'h6019: out_word = 8'hCD;
		16'h601A: out_word = 8'hB1;
		16'h601B: out_word = 8'h20;
		16'h601C: out_word = 8'h16;
		16'h601D: out_word = 8'hFE;
		16'h601E: out_word = 8'hCD;
		16'h601F: out_word = 8'hAF;
		16'h6020: out_word = 8'h20;
		16'h6021: out_word = 8'h53;
		16'h6022: out_word = 8'hCD;
		16'h6023: out_word = 8'hAF;
		16'h6024: out_word = 8'h20;
		16'h6025: out_word = 8'h16;
		16'h6026: out_word = 8'h00;
		16'h6027: out_word = 8'hCD;
		16'h6028: out_word = 8'hAF;
		16'h6029: out_word = 8'h20;
		16'h602A: out_word = 8'h56;
		16'h602B: out_word = 8'hCD;
		16'h602C: out_word = 8'hAF;
		16'h602D: out_word = 8'h20;
		16'h602E: out_word = 8'h16;
		16'h602F: out_word = 8'h01;
		16'h6030: out_word = 8'hCD;
		16'h6031: out_word = 8'hAF;
		16'h6032: out_word = 8'h20;
		16'h6033: out_word = 8'h16;
		16'h6034: out_word = 8'hF7;
		16'h6035: out_word = 8'hCD;
		16'h6036: out_word = 8'hAF;
		16'h6037: out_word = 8'h20;
		16'h6038: out_word = 8'h06;
		16'h6039: out_word = 8'h16;
		16'h603A: out_word = 8'h16;
		16'h603B: out_word = 8'h4E;
		16'h603C: out_word = 8'hCD;
		16'h603D: out_word = 8'hB1;
		16'h603E: out_word = 8'h20;
		16'h603F: out_word = 8'h06;
		16'h6040: out_word = 8'h0C;
		16'h6041: out_word = 8'h16;
		16'h6042: out_word = 8'h00;
		16'h6043: out_word = 8'hCD;
		16'h6044: out_word = 8'hB1;
		16'h6045: out_word = 8'h20;
		16'h6046: out_word = 8'h06;
		16'h6047: out_word = 8'h03;
		16'h6048: out_word = 8'h16;
		16'h6049: out_word = 8'hF5;
		16'h604A: out_word = 8'hCD;
		16'h604B: out_word = 8'hB1;
		16'h604C: out_word = 8'h20;
		16'h604D: out_word = 8'h16;
		16'h604E: out_word = 8'hFB;
		16'h604F: out_word = 8'hCD;
		16'h6050: out_word = 8'hAF;
		16'h6051: out_word = 8'h20;
		16'h6052: out_word = 8'h06;
		16'h6053: out_word = 8'h00;
		16'h6054: out_word = 8'h16;
		16'h6055: out_word = 8'h00;
		16'h6056: out_word = 8'hCD;
		16'h6057: out_word = 8'hB1;
		16'h6058: out_word = 8'h20;
		16'h6059: out_word = 8'h16;
		16'h605A: out_word = 8'hF7;
		16'h605B: out_word = 8'hCD;
		16'h605C: out_word = 8'hAF;
		16'h605D: out_word = 8'h20;
		16'h605E: out_word = 8'h06;
		16'h605F: out_word = 8'h32;
		16'h6060: out_word = 8'h16;
		16'h6061: out_word = 8'h4E;
		16'h6062: out_word = 8'hCD;
		16'h6063: out_word = 8'hB1;
		16'h6064: out_word = 8'h20;
		16'h6065: out_word = 8'h7E;
		16'h6066: out_word = 8'h23;
		16'h6067: out_word = 8'hFE;
		16'h6068: out_word = 8'h10;
		16'h6069: out_word = 8'h20;
		16'h606A: out_word = 8'h9C;
		16'h606B: out_word = 8'h06;
		16'h606C: out_word = 8'h00;
		16'h606D: out_word = 8'hCD;
		16'h606E: out_word = 8'hB1;
		16'h606F: out_word = 8'h20;
		16'h6070: out_word = 8'hFA;
		16'h6071: out_word = 8'h76;
		16'h6072: out_word = 8'h20;
		16'h6073: out_word = 8'hCD;
		16'h6074: out_word = 8'hB1;
		16'h6075: out_word = 8'h20;
		16'h6076: out_word = 8'hDB;
		16'h6077: out_word = 8'h1F;
		16'h6078: out_word = 8'hE6;
		16'h6079: out_word = 8'h40;
		16'h607A: out_word = 8'hC2;
		16'h607B: out_word = 8'h39;
		16'h607C: out_word = 8'h3F;
		16'h607D: out_word = 8'h3A;
		16'h607E: out_word = 8'hD8;
		16'h607F: out_word = 8'h5C;
		16'h6080: out_word = 8'hB7;
		16'h6081: out_word = 8'hC0;
		16'h6082: out_word = 8'h0E;
		16'h6083: out_word = 8'h7F;
		16'h6084: out_word = 8'h7B;
		16'h6085: out_word = 8'hD3;
		16'h6086: out_word = 8'h3F;
		16'h6087: out_word = 8'hCD;
		16'h6088: out_word = 8'hBE;
		16'h6089: out_word = 8'h33;
		16'h608A: out_word = 8'h06;
		16'h608B: out_word = 8'h03;
		16'h608C: out_word = 8'h7E;
		16'h608D: out_word = 8'hD3;
		16'h608E: out_word = 8'h5F;
		16'h608F: out_word = 8'hE5;
		16'h6090: out_word = 8'hF3;
		16'h6091: out_word = 8'h3E;
		16'h6092: out_word = 8'h80;
		16'h6093: out_word = 8'hD3;
		16'h6094: out_word = 8'h1F;
		16'h6095: out_word = 8'hC5;
		16'h6096: out_word = 8'hCD;
		16'h6097: out_word = 8'hE5;
		16'h6098: out_word = 8'h3F;
		16'h6099: out_word = 8'hDB;
		16'h609A: out_word = 8'h1F;
		16'h609B: out_word = 8'hE6;
		16'h609C: out_word = 8'h7F;
		16'h609D: out_word = 8'hC1;
		16'h609E: out_word = 8'h28;
		16'h609F: out_word = 8'h06;
		16'h60A0: out_word = 8'h10;
		16'h60A1: out_word = 8'hEE;
		16'h60A2: out_word = 8'h21;
		16'h60A3: out_word = 8'hD6;
		16'h60A4: out_word = 8'h5C;
		16'h60A5: out_word = 8'h34;
		16'h60A6: out_word = 8'hE1;
		16'h60A7: out_word = 8'h7E;
		16'h60A8: out_word = 8'h23;
		16'h60A9: out_word = 8'hFE;
		16'h60AA: out_word = 8'h01;
		16'h60AB: out_word = 8'h20;
		16'h60AC: out_word = 8'hDD;
		16'h60AD: out_word = 8'hFB;
		16'h60AE: out_word = 8'hC9;
		16'h60AF: out_word = 8'h06;
		16'h60B0: out_word = 8'h01;
		16'h60B1: out_word = 8'hDB;
		16'h60B2: out_word = 8'hFF;
		16'h60B3: out_word = 8'hE6;
		16'h60B4: out_word = 8'hC0;
		16'h60B5: out_word = 8'h28;
		16'h60B6: out_word = 8'hFA;
		16'h60B7: out_word = 8'hF8;
		16'h60B8: out_word = 8'hED;
		16'h60B9: out_word = 8'h51;
		16'h60BA: out_word = 8'h10;
		16'h60BB: out_word = 8'hF5;
		16'h60BC: out_word = 8'hC9;
		16'h60BD: out_word = 8'h21;
		16'h60BE: out_word = 8'hD7;
		16'h60BF: out_word = 8'h5C;
		16'h60C0: out_word = 8'h46;
		16'h60C1: out_word = 8'hCD;
		16'h60C2: out_word = 8'hEA;
		16'h60C3: out_word = 8'h32;
		16'h60C4: out_word = 8'h1E;
		16'h60C5: out_word = 8'hFF;
		16'h60C6: out_word = 8'hC5;
		16'h60C7: out_word = 8'h1C;
		16'h60C8: out_word = 8'h7B;
		16'h60C9: out_word = 8'h06;
		16'h60CA: out_word = 8'h1B;
		16'h60CB: out_word = 8'hCD;
		16'h60CC: out_word = 8'h24;
		16'h60CD: out_word = 8'h32;
		16'h60CE: out_word = 8'hCD;
		16'h60CF: out_word = 8'hEB;
		16'h60D0: out_word = 8'h1F;
		16'h60D1: out_word = 8'hCD;
		16'h60D2: out_word = 8'hF6;
		16'h60D3: out_word = 8'h32;
		16'h60D4: out_word = 8'h3A;
		16'h60D5: out_word = 8'hDA;
		16'h60D6: out_word = 8'h5C;
		16'h60D7: out_word = 8'hFE;
		16'h60D8: out_word = 8'h80;
		16'h60D9: out_word = 8'h20;
		16'h60DA: out_word = 8'h06;
		16'h60DB: out_word = 8'hCD;
		16'h60DC: out_word = 8'hF6;
		16'h60DD: out_word = 8'h1F;
		16'h60DE: out_word = 8'hCD;
		16'h60DF: out_word = 8'hF1;
		16'h60E0: out_word = 8'h32;
		16'h60E1: out_word = 8'hC1;
		16'h60E2: out_word = 8'h10;
		16'h60E3: out_word = 8'hE2;
		16'h60E4: out_word = 8'hC9;
		16'h60E5: out_word = 8'hF5;
		16'h60E6: out_word = 8'h3A;
		16'h60E7: out_word = 8'hF8;
		16'h60E8: out_word = 8'h5C;
		16'h60E9: out_word = 8'hFE;
		16'h60EA: out_word = 8'hFF;
		16'h60EB: out_word = 8'h28;
		16'h60EC: out_word = 8'h2F;
		16'h60ED: out_word = 8'hF1;
		16'h60EE: out_word = 8'hCD;
		16'h60EF: out_word = 8'h70;
		16'h60F0: out_word = 8'h29;
		16'h60F1: out_word = 8'hF5;
		16'h60F2: out_word = 8'h3A;
		16'h60F3: out_word = 8'hB6;
		16'h60F4: out_word = 8'h5C;
		16'h60F5: out_word = 8'hFE;
		16'h60F6: out_word = 8'hF4;
		16'h60F7: out_word = 8'h28;
		16'h60F8: out_word = 8'h23;
		16'h60F9: out_word = 8'hAF;
		16'h60FA: out_word = 8'h21;
		16'h60FB: out_word = 8'h18;
		16'h60FC: out_word = 8'h5D;
		16'h60FD: out_word = 8'hB6;
		16'h60FE: out_word = 8'h36;
		16'h60FF: out_word = 8'hFF;
		16'h6100: out_word = 8'h28;
		16'h6101: out_word = 8'h1A;
		16'h6102: out_word = 8'h3A;
		16'h6103: out_word = 8'h0C;
		16'h6104: out_word = 8'h5D;
		16'h6105: out_word = 8'hB7;
		16'h6106: out_word = 8'h21;
		16'h6107: out_word = 8'hC3;
		16'h6108: out_word = 8'h5C;
		16'h6109: out_word = 8'h11;
		16'h610A: out_word = 8'h33;
		16'h610B: out_word = 8'h5D;
		16'h610C: out_word = 8'h20;
		16'h610D: out_word = 8'h03;
		16'h610E: out_word = 8'h11;
		16'h610F: out_word = 8'h34;
		16'h6110: out_word = 8'h5E;
		16'h6111: out_word = 8'h06;
		16'h6112: out_word = 8'h2D;
		16'h6113: out_word = 8'h4E;
		16'h6114: out_word = 8'h1A;
		16'h6115: out_word = 8'h77;
		16'h6116: out_word = 8'h79;
		16'h6117: out_word = 8'h12;
		16'h6118: out_word = 8'h23;
		16'h6119: out_word = 8'h13;
		16'h611A: out_word = 8'h10;
		16'h611B: out_word = 8'hF7;
		16'h611C: out_word = 8'hF1;
		16'h611D: out_word = 8'hC9;
		16'h611E: out_word = 8'h2A;
		16'h611F: out_word = 8'h59;
		16'h6120: out_word = 8'h5C;
		16'h6121: out_word = 8'h36;
		16'h6122: out_word = 8'h0D;
		16'h6123: out_word = 8'h22;
		16'h6124: out_word = 8'h5B;
		16'h6125: out_word = 8'h5C;
		16'h6126: out_word = 8'h23;
		16'h6127: out_word = 8'h36;
		16'h6128: out_word = 8'h80;
		16'h6129: out_word = 8'hC9;
		16'h612A: out_word = 8'hED;
		16'h612B: out_word = 8'h5B;
		16'h612C: out_word = 8'h59;
		16'h612D: out_word = 8'h5C;
		16'h612E: out_word = 8'h21;
		16'h612F: out_word = 8'h20;
		16'h6130: out_word = 8'h5D;
		16'h6131: out_word = 8'hCD;
		16'h6132: out_word = 8'hB0;
		16'h6133: out_word = 8'h02;
		16'h6134: out_word = 8'hC9;
		16'h6135: out_word = 8'h3A;
		16'h6136: out_word = 8'h0F;
		16'h6137: out_word = 8'h5D;
		16'h6138: out_word = 8'hB7;
		16'h6139: out_word = 8'hF5;
		16'h613A: out_word = 8'hC4;
		16'h613B: out_word = 8'h2A;
		16'h613C: out_word = 8'h21;
		16'h613D: out_word = 8'hF1;
		16'h613E: out_word = 8'hCC;
		16'h613F: out_word = 8'h1E;
		16'h6140: out_word = 8'h21;
		16'h6141: out_word = 8'h2A;
		16'h6142: out_word = 8'h59;
		16'h6143: out_word = 8'h5C;
		16'h6144: out_word = 8'hCD;
		16'h6145: out_word = 8'h80;
		16'h6146: out_word = 8'h3D;
		16'h6147: out_word = 8'h3A;
		16'h6148: out_word = 8'h19;
		16'h6149: out_word = 8'h5D;
		16'h614A: out_word = 8'hC6;
		16'h614B: out_word = 8'h41;
		16'h614C: out_word = 8'hD7;
		16'h614D: out_word = 8'h3E;
		16'h614E: out_word = 8'h3E;
		16'h614F: out_word = 8'hD7;
		16'h6150: out_word = 8'hFD;
		16'h6151: out_word = 8'h36;
		16'h6152: out_word = 8'h00;
		16'h6153: out_word = 8'hFF;
		16'h6154: out_word = 8'hFB;
		16'h6155: out_word = 8'hC3;
		16'h6156: out_word = 8'h80;
		16'h6157: out_word = 8'h3B;
		16'h6158: out_word = 8'hCD;
		16'h6159: out_word = 8'h2A;
		16'h615A: out_word = 8'h1E;
		16'h615B: out_word = 8'hCD;
		16'h615C: out_word = 8'h8C;
		16'h615D: out_word = 8'h1D;
		16'h615E: out_word = 8'hFE;
		16'h615F: out_word = 8'h2C;
		16'h6160: out_word = 8'hC2;
		16'h6161: out_word = 8'h1A;
		16'h6162: out_word = 8'h1D;
		16'h6163: out_word = 8'h2A;
		16'h6164: out_word = 8'hDB;
		16'h6165: out_word = 8'h5C;
		16'h6166: out_word = 8'h22;
		16'h6167: out_word = 8'hD9;
		16'h6168: out_word = 8'h5C;
		16'h6169: out_word = 8'hCD;
		16'h616A: out_word = 8'h0B;
		16'h616B: out_word = 8'h1E;
		16'h616C: out_word = 8'hCD;
		16'h616D: out_word = 8'h75;
		16'h616E: out_word = 8'h1D;
		16'h616F: out_word = 8'h2A;
		16'h6170: out_word = 8'hDB;
		16'h6171: out_word = 8'h5C;
		16'h6172: out_word = 8'h7C;
		16'h6173: out_word = 8'hB7;
		16'h6174: out_word = 8'hC2;
		16'h6175: out_word = 8'h1A;
		16'h6176: out_word = 8'h1D;
		16'h6177: out_word = 8'h23;
		16'h6178: out_word = 8'h22;
		16'h6179: out_word = 8'hD7;
		16'h617A: out_word = 8'h5C;
		16'h617B: out_word = 8'h2A;
		16'h617C: out_word = 8'hD9;
		16'h617D: out_word = 8'h5C;
		16'h617E: out_word = 8'h22;
		16'h617F: out_word = 8'hDB;
		16'h6180: out_word = 8'h5C;
		16'h6181: out_word = 8'hC9;
		16'h6182: out_word = 8'h2A;
		16'h6183: out_word = 8'h11;
		16'h6184: out_word = 8'h5D;
		16'h6185: out_word = 8'h22;
		16'h6186: out_word = 8'h5D;
		16'h6187: out_word = 8'h5C;
		16'h6188: out_word = 8'hCD;
		16'h6189: out_word = 8'h0B;
		16'h618A: out_word = 8'h1E;
		16'h618B: out_word = 8'hCD;
		16'h618C: out_word = 8'hD0;
		16'h618D: out_word = 8'h1D;
		16'h618E: out_word = 8'hCD;
		16'h618F: out_word = 8'h8C;
		16'h6190: out_word = 8'h1D;
		16'h6191: out_word = 8'hFE;
		16'h6192: out_word = 8'h41;
		16'h6193: out_word = 8'h30;
		16'h6194: out_word = 8'h05;
		16'h6195: out_word = 8'hCD;
		16'h6196: out_word = 8'h2A;
		16'h6197: out_word = 8'h1E;
		16'h6198: out_word = 8'h18;
		16'h6199: out_word = 8'hF4;
		16'h619A: out_word = 8'hFE;
		16'h619B: out_word = 8'hA5;
		16'h619C: out_word = 8'hF5;
		16'h619D: out_word = 8'hCC;
		16'h619E: out_word = 8'h58;
		16'h619F: out_word = 8'h21;
		16'h61A0: out_word = 8'hF1;
		16'h61A1: out_word = 8'h28;
		16'h61A2: out_word = 8'h0B;
		16'h61A3: out_word = 8'hE6;
		16'h61A4: out_word = 8'hDF;
		16'h61A5: out_word = 8'hFE;
		16'h61A6: out_word = 8'h52;
		16'h61A7: out_word = 8'h28;
		16'h61A8: out_word = 8'h05;
		16'h61A9: out_word = 8'hFE;
		16'h61AA: out_word = 8'h57;
		16'h61AB: out_word = 8'hC2;
		16'h61AC: out_word = 8'h1A;
		16'h61AD: out_word = 8'h1D;
		16'h61AE: out_word = 8'h32;
		16'h61AF: out_word = 8'h09;
		16'h61B0: out_word = 8'h5D;
		16'h61B1: out_word = 8'hCD;
		16'h61B2: out_word = 8'h75;
		16'h61B3: out_word = 8'h1D;
		16'h61B4: out_word = 8'h3E;
		16'h61B5: out_word = 8'h23;
		16'h61B6: out_word = 8'h32;
		16'h61B7: out_word = 8'hE5;
		16'h61B8: out_word = 8'h5C;
		16'h61B9: out_word = 8'h3E;
		16'h61BA: out_word = 8'h00;
		16'h61BB: out_word = 8'h32;
		16'h61BC: out_word = 8'hE6;
		16'h61BD: out_word = 8'h5C;
		16'h61BE: out_word = 8'hCD;
		16'h61BF: out_word = 8'hDB;
		16'h61C0: out_word = 8'h21;
		16'h61C1: out_word = 8'hF5;
		16'h61C2: out_word = 8'hCD;
		16'h61C3: out_word = 8'h0F;
		16'h61C4: out_word = 8'h22;
		16'h61C5: out_word = 8'hF1;
		16'h61C6: out_word = 8'hF5;
		16'h61C7: out_word = 8'hC4;
		16'h61C8: out_word = 8'h88;
		16'h61C9: out_word = 8'h22;
		16'h61CA: out_word = 8'hF1;
		16'h61CB: out_word = 8'hCD;
		16'h61CC: out_word = 8'h42;
		16'h61CD: out_word = 8'h22;
		16'h61CE: out_word = 8'h2A;
		16'h61CF: out_word = 8'h11;
		16'h61D0: out_word = 8'h5D;
		16'h61D1: out_word = 8'h01;
		16'h61D2: out_word = 8'h24;
		16'h61D3: out_word = 8'h01;
		16'h61D4: out_word = 8'h09;
		16'h61D5: out_word = 8'h22;
		16'h61D6: out_word = 8'h11;
		16'h61D7: out_word = 8'h5D;
		16'h61D8: out_word = 8'hC3;
		16'h61D9: out_word = 8'hD3;
		16'h61DA: out_word = 8'h01;
		16'h61DB: out_word = 8'h3E;
		16'h61DC: out_word = 8'h0A;
		16'h61DD: out_word = 8'h32;
		16'h61DE: out_word = 8'h06;
		16'h61DF: out_word = 8'h5D;
		16'h61E0: out_word = 8'hCD;
		16'h61E1: out_word = 8'hB0;
		16'h61E2: out_word = 8'h1C;
		16'h61E3: out_word = 8'hF5;
		16'h61E4: out_word = 8'hCD;
		16'h61E5: out_word = 8'h05;
		16'h61E6: out_word = 8'h04;
		16'h61E7: out_word = 8'hF1;
		16'h61E8: out_word = 8'h20;
		16'h61E9: out_word = 8'h1C;
		16'h61EA: out_word = 8'h3A;
		16'h61EB: out_word = 8'h09;
		16'h61EC: out_word = 8'h5D;
		16'h61ED: out_word = 8'hFE;
		16'h61EE: out_word = 8'h52;
		16'h61EF: out_word = 8'h28;
		16'h61F0: out_word = 8'h10;
		16'h61F1: out_word = 8'h21;
		16'h61F2: out_word = 8'hE6;
		16'h61F3: out_word = 8'h5C;
		16'h61F4: out_word = 8'h34;
		16'h61F5: out_word = 8'hCD;
		16'h61F6: out_word = 8'hB3;
		16'h61F7: out_word = 8'h1C;
		16'h61F8: out_word = 8'h28;
		16'h61F9: out_word = 8'hF7;
		16'h61FA: out_word = 8'h21;
		16'h61FB: out_word = 8'hE6;
		16'h61FC: out_word = 8'h5C;
		16'h61FD: out_word = 8'h35;
		16'h61FE: out_word = 8'hCD;
		16'h61FF: out_word = 8'hB3;
		16'h6200: out_word = 8'h1C;
		16'h6201: out_word = 8'hCD;
		16'h6202: out_word = 8'h5D;
		16'h6203: out_word = 8'h16;
		16'h6204: out_word = 8'hAF;
		16'h6205: out_word = 8'hC9;
		16'h6206: out_word = 8'h3A;
		16'h6207: out_word = 8'h09;
		16'h6208: out_word = 8'h5D;
		16'h6209: out_word = 8'hFE;
		16'h620A: out_word = 8'h52;
		16'h620B: out_word = 8'hC0;
		16'h620C: out_word = 8'hC3;
		16'h620D: out_word = 8'hD9;
		16'h620E: out_word = 8'h03;
		16'h620F: out_word = 8'h3A;
		16'h6210: out_word = 8'hDB;
		16'h6211: out_word = 8'h5C;
		16'h6212: out_word = 8'hE7;
		16'h6213: out_word = 8'h27;
		16'h6214: out_word = 8'h17;
		16'h6215: out_word = 8'h78;
		16'h6216: out_word = 8'hB1;
		16'h6217: out_word = 8'hC2;
		16'h6218: out_word = 8'h1B;
		16'h6219: out_word = 8'h22;
		16'h621A: out_word = 8'hC9;
		16'h621B: out_word = 8'h3E;
		16'h621C: out_word = 8'h19;
		16'h621D: out_word = 8'h32;
		16'h621E: out_word = 8'h3A;
		16'h621F: out_word = 8'h5C;
		16'h6220: out_word = 8'h21;
		16'h6221: out_word = 8'h04;
		16'h6222: out_word = 8'h28;
		16'h6223: out_word = 8'h3E;
		16'h6224: out_word = 8'h0A;
		16'h6225: out_word = 8'hC3;
		16'h6226: out_word = 8'h4A;
		16'h6227: out_word = 8'h1C;
		16'h6228: out_word = 8'h3E;
		16'h6229: out_word = 8'h0B;
		16'h622A: out_word = 8'h21;
		16'h622B: out_word = 8'h12;
		16'h622C: out_word = 8'h28;
		16'h622D: out_word = 8'h18;
		16'h622E: out_word = 8'hF6;
		16'h622F: out_word = 8'hE5;
		16'h6230: out_word = 8'h0E;
		16'h6231: out_word = 8'h20;
		16'h6232: out_word = 8'hEF;
		16'h6233: out_word = 8'h3A;
		16'h6234: out_word = 8'hD7;
		16'h6235: out_word = 8'h5C;
		16'h6236: out_word = 8'h77;
		16'h6237: out_word = 8'h23;
		16'h6238: out_word = 8'hAF;
		16'h6239: out_word = 8'h77;
		16'h623A: out_word = 8'h23;
		16'h623B: out_word = 8'h77;
		16'h623C: out_word = 8'h23;
		16'h623D: out_word = 8'h77;
		16'h623E: out_word = 8'h3E;
		16'h623F: out_word = 8'h7F;
		16'h6240: out_word = 8'hE1;
		16'h6241: out_word = 8'hC9;
		16'h6242: out_word = 8'hF5;
		16'h6243: out_word = 8'hCD;
		16'h6244: out_word = 8'h0F;
		16'h6245: out_word = 8'h22;
		16'h6246: out_word = 8'hEB;
		16'h6247: out_word = 8'h2A;
		16'h6248: out_word = 8'h53;
		16'h6249: out_word = 8'h5C;
		16'h624A: out_word = 8'hED;
		16'h624B: out_word = 8'h4B;
		16'h624C: out_word = 8'h4F;
		16'h624D: out_word = 8'h5C;
		16'h624E: out_word = 8'hED;
		16'h624F: out_word = 8'h42;
		16'h6250: out_word = 8'hEB;
		16'h6251: out_word = 8'h73;
		16'h6252: out_word = 8'h23;
		16'h6253: out_word = 8'h72;
		16'h6254: out_word = 8'hCD;
		16'h6255: out_word = 8'hB2;
		16'h6256: out_word = 8'h22;
		16'h6257: out_word = 8'h3A;
		16'h6258: out_word = 8'h09;
		16'h6259: out_word = 8'h5D;
		16'h625A: out_word = 8'hFE;
		16'h625B: out_word = 8'hA5;
		16'h625C: out_word = 8'hCC;
		16'h625D: out_word = 8'h2F;
		16'h625E: out_word = 8'h22;
		16'h625F: out_word = 8'h28;
		16'h6260: out_word = 8'h0A;
		16'h6261: out_word = 8'h3A;
		16'h6262: out_word = 8'h09;
		16'h6263: out_word = 8'h5D;
		16'h6264: out_word = 8'hFE;
		16'h6265: out_word = 8'h52;
		16'h6266: out_word = 8'h3E;
		16'h6267: out_word = 8'hFF;
		16'h6268: out_word = 8'h20;
		16'h6269: out_word = 8'h01;
		16'h626A: out_word = 8'hAF;
		16'h626B: out_word = 8'h77;
		16'h626C: out_word = 8'hF1;
		16'h626D: out_word = 8'hC3;
		16'h626E: out_word = 8'h70;
		16'h626F: out_word = 8'h22;
		16'h6270: out_word = 8'hF5;
		16'h6271: out_word = 8'h01;
		16'h6272: out_word = 8'h14;
		16'h6273: out_word = 8'h00;
		16'h6274: out_word = 8'h09;
		16'h6275: out_word = 8'hE5;
		16'h6276: out_word = 8'hCD;
		16'h6277: out_word = 8'h23;
		16'h6278: out_word = 8'h24;
		16'h6279: out_word = 8'hE1;
		16'h627A: out_word = 8'h23;
		16'h627B: out_word = 8'h06;
		16'h627C: out_word = 8'h01;
		16'h627D: out_word = 8'hF1;
		16'h627E: out_word = 8'hB7;
		16'h627F: out_word = 8'hF5;
		16'h6280: out_word = 8'hC4;
		16'h6281: out_word = 8'h4D;
		16'h6282: out_word = 8'h1E;
		16'h6283: out_word = 8'hF1;
		16'h6284: out_word = 8'hCC;
		16'h6285: out_word = 8'h3D;
		16'h6286: out_word = 8'h1E;
		16'h6287: out_word = 8'hC9;
		16'h6288: out_word = 8'h2A;
		16'h6289: out_word = 8'hD7;
		16'h628A: out_word = 8'h5C;
		16'h628B: out_word = 8'hE5;
		16'h628C: out_word = 8'h21;
		16'h628D: out_word = 8'h00;
		16'h628E: out_word = 8'h20;
		16'h628F: out_word = 8'h22;
		16'h6290: out_word = 8'hD7;
		16'h6291: out_word = 8'h5C;
		16'h6292: out_word = 8'hCD;
		16'h6293: out_word = 8'h9A;
		16'h6294: out_word = 8'h22;
		16'h6295: out_word = 8'hE1;
		16'h6296: out_word = 8'h22;
		16'h6297: out_word = 8'hD7;
		16'h6298: out_word = 8'h5C;
		16'h6299: out_word = 8'hC9;
		16'h629A: out_word = 8'h21;
		16'h629B: out_word = 8'h00;
		16'h629C: out_word = 8'h10;
		16'h629D: out_word = 8'h22;
		16'h629E: out_word = 8'hD9;
		16'h629F: out_word = 8'h5C;
		16'h62A0: out_word = 8'hCD;
		16'h62A1: out_word = 8'hC4;
		16'h62A2: out_word = 8'h1A;
		16'h62A3: out_word = 8'hCD;
		16'h62A4: out_word = 8'h59;
		16'h62A5: out_word = 8'h1B;
		16'h62A6: out_word = 8'h21;
		16'h62A7: out_word = 8'h00;
		16'h62A8: out_word = 8'h00;
		16'h62A9: out_word = 8'h22;
		16'h62AA: out_word = 8'hE8;
		16'h62AB: out_word = 8'h5C;
		16'h62AC: out_word = 8'hCD;
		16'h62AD: out_word = 8'h6B;
		16'h62AE: out_word = 8'h16;
		16'h62AF: out_word = 8'hC3;
		16'h62B0: out_word = 8'h43;
		16'h62B1: out_word = 8'h1E;
		16'h62B2: out_word = 8'h2A;
		16'h62B3: out_word = 8'h53;
		16'h62B4: out_word = 8'h5C;
		16'h62B5: out_word = 8'h2B;
		16'h62B6: out_word = 8'h22;
		16'h62B7: out_word = 8'h51;
		16'h62B8: out_word = 8'h5C;
		16'h62B9: out_word = 8'hE5;
		16'h62BA: out_word = 8'h01;
		16'h62BB: out_word = 8'h24;
		16'h62BC: out_word = 8'h01;
		16'h62BD: out_word = 8'hCD;
		16'h62BE: out_word = 8'h32;
		16'h62BF: out_word = 8'h1E;
		16'h62C0: out_word = 8'h3E;
		16'h62C1: out_word = 8'h00;
		16'h62C2: out_word = 8'h06;
		16'h62C3: out_word = 8'h00;
		16'h62C4: out_word = 8'h12;
		16'h62C5: out_word = 8'h1B;
		16'h62C6: out_word = 8'h10;
		16'h62C7: out_word = 8'hFC;
		16'h62C8: out_word = 8'hE1;
		16'h62C9: out_word = 8'hE5;
		16'h62CA: out_word = 8'h11;
		16'h62CB: out_word = 8'h0E;
		16'h62CC: out_word = 8'h3D;
		16'h62CD: out_word = 8'h73;
		16'h62CE: out_word = 8'h23;
		16'h62CF: out_word = 8'h72;
		16'h62D0: out_word = 8'h23;
		16'h62D1: out_word = 8'h11;
		16'h62D2: out_word = 8'h06;
		16'h62D3: out_word = 8'h3D;
		16'h62D4: out_word = 8'h73;
		16'h62D5: out_word = 8'h23;
		16'h62D6: out_word = 8'h72;
		16'h62D7: out_word = 8'h23;
		16'h62D8: out_word = 8'h36;
		16'h62D9: out_word = 8'h44;
		16'h62DA: out_word = 8'h23;
		16'h62DB: out_word = 8'h23;
		16'h62DC: out_word = 8'h23;
		16'h62DD: out_word = 8'h23;
		16'h62DE: out_word = 8'h23;
		16'h62DF: out_word = 8'h36;
		16'h62E0: out_word = 8'h24;
		16'h62E1: out_word = 8'h23;
		16'h62E2: out_word = 8'h36;
		16'h62E3: out_word = 8'h01;
		16'h62E4: out_word = 8'h23;
		16'h62E5: out_word = 8'h3A;
		16'h62E6: out_word = 8'hF6;
		16'h62E7: out_word = 8'h5C;
		16'h62E8: out_word = 8'h77;
		16'h62E9: out_word = 8'h23;
		16'h62EA: out_word = 8'h3A;
		16'h62EB: out_word = 8'h1E;
		16'h62EC: out_word = 8'h5D;
		16'h62ED: out_word = 8'h77;
		16'h62EE: out_word = 8'h23;
		16'h62EF: out_word = 8'h3A;
		16'h62F0: out_word = 8'h09;
		16'h62F1: out_word = 8'h5D;
		16'h62F2: out_word = 8'hFE;
		16'h62F3: out_word = 8'h52;
		16'h62F4: out_word = 8'h36;
		16'h62F5: out_word = 8'h00;
		16'h62F6: out_word = 8'h28;
		16'h62F7: out_word = 8'h04;
		16'h62F8: out_word = 8'h3A;
		16'h62F9: out_word = 8'hE8;
		16'h62FA: out_word = 8'h5C;
		16'h62FB: out_word = 8'h77;
		16'h62FC: out_word = 8'h23;
		16'h62FD: out_word = 8'h70;
		16'h62FE: out_word = 8'h28;
		16'h62FF: out_word = 8'h04;
		16'h6300: out_word = 8'h3A;
		16'h6301: out_word = 8'hE9;
		16'h6302: out_word = 8'h5C;
		16'h6303: out_word = 8'h77;
		16'h6304: out_word = 8'h23;
		16'h6305: out_word = 8'hEB;
		16'h6306: out_word = 8'hE1;
		16'h6307: out_word = 8'hD5;
		16'h6308: out_word = 8'h11;
		16'h6309: out_word = 8'h10;
		16'h630A: out_word = 8'h00;
		16'h630B: out_word = 8'h19;
		16'h630C: out_word = 8'hEB;
		16'h630D: out_word = 8'h21;
		16'h630E: out_word = 8'hDD;
		16'h630F: out_word = 8'h5C;
		16'h6310: out_word = 8'h01;
		16'h6311: out_word = 8'h10;
		16'h6312: out_word = 8'h00;
		16'h6313: out_word = 8'hED;
		16'h6314: out_word = 8'hB0;
		16'h6315: out_word = 8'hE1;
		16'h6316: out_word = 8'hC9;
		16'h6317: out_word = 8'h0E;
		16'h6318: out_word = 8'h0D;
		16'h6319: out_word = 8'hEF;
		16'h631A: out_word = 8'h4E;
		16'h631B: out_word = 8'hEF;
		16'h631C: out_word = 8'h01;
		16'h631D: out_word = 8'h24;
		16'h631E: out_word = 8'h00;
		16'h631F: out_word = 8'h09;
		16'h6320: out_word = 8'hC9;
		16'h6321: out_word = 8'h0E;
		16'h6322: out_word = 8'h24;
		16'h6323: out_word = 8'h06;
		16'h6324: out_word = 8'h00;
		16'h6325: out_word = 8'h2A;
		16'h6326: out_word = 8'h51;
		16'h6327: out_word = 8'h5C;
		16'h6328: out_word = 8'h09;
		16'h6329: out_word = 8'hC9;
		16'h632A: out_word = 8'h0E;
		16'h632B: out_word = 8'h0D;
		16'h632C: out_word = 8'hEF;
		16'h632D: out_word = 8'h34;
		16'h632E: out_word = 8'hC0;
		16'h632F: out_word = 8'hE5;
		16'h6330: out_word = 8'hCD;
		16'h6331: out_word = 8'h43;
		16'h6332: out_word = 8'h24;
		16'h6333: out_word = 8'hCD;
		16'h6334: out_word = 8'hFC;
		16'h6335: out_word = 8'h23;
		16'h6336: out_word = 8'hE1;
		16'h6337: out_word = 8'h23;
		16'h6338: out_word = 8'h34;
		16'h6339: out_word = 8'hE5;
		16'h633A: out_word = 8'hCD;
		16'h633B: out_word = 8'h18;
		16'h633C: out_word = 8'h24;
		16'h633D: out_word = 8'hE1;
		16'h633E: out_word = 8'h3E;
		16'h633F: out_word = 8'h10;
		16'h6340: out_word = 8'hBE;
		16'h6341: out_word = 8'hC0;
		16'h6342: out_word = 8'hE5;
		16'h6343: out_word = 8'h0E;
		16'h6344: out_word = 8'h0F;
		16'h6345: out_word = 8'hEF;
		16'h6346: out_word = 8'h7E;
		16'h6347: out_word = 8'hFE;
		16'h6348: out_word = 8'h7F;
		16'h6349: out_word = 8'hE1;
		16'h634A: out_word = 8'h28;
		16'h634B: out_word = 8'h0C;
		16'h634C: out_word = 8'h2A;
		16'h634D: out_word = 8'h51;
		16'h634E: out_word = 8'h5C;
		16'h634F: out_word = 8'hCD;
		16'h6350: out_word = 8'hE1;
		16'h6351: out_word = 8'h26;
		16'h6352: out_word = 8'h0E;
		16'h6353: out_word = 8'h0E;
		16'h6354: out_word = 8'hEF;
		16'h6355: out_word = 8'hC3;
		16'h6356: out_word = 8'h79;
		16'h6357: out_word = 8'h23;
		16'h6358: out_word = 8'hCD;
		16'h6359: out_word = 8'hCF;
		16'h635A: out_word = 8'h23;
		16'h635B: out_word = 8'hF5;
		16'h635C: out_word = 8'hCC;
		16'h635D: out_word = 8'h18;
		16'h635E: out_word = 8'h24;
		16'h635F: out_word = 8'h0E;
		16'h6360: out_word = 8'h0E;
		16'h6361: out_word = 8'hEF;
		16'h6362: out_word = 8'hF1;
		16'h6363: out_word = 8'hC4;
		16'h6364: out_word = 8'h70;
		16'h6365: out_word = 8'h23;
		16'h6366: out_word = 8'hC9;
		16'h6367: out_word = 8'h36;
		16'h6368: out_word = 8'h00;
		16'h6369: out_word = 8'h0E;
		16'h636A: out_word = 8'h19;
		16'h636B: out_word = 8'hEF;
		16'h636C: out_word = 8'h16;
		16'h636D: out_word = 8'h20;
		16'h636E: out_word = 8'h5E;
		16'h636F: out_word = 8'hC9;
		16'h6370: out_word = 8'hCD;
		16'h6371: out_word = 8'h67;
		16'h6372: out_word = 8'h23;
		16'h6373: out_word = 8'hED;
		16'h6374: out_word = 8'h53;
		16'h6375: out_word = 8'hD7;
		16'h6376: out_word = 8'h5C;
		16'h6377: out_word = 8'h18;
		16'h6378: out_word = 8'h08;
		16'h6379: out_word = 8'hCD;
		16'h637A: out_word = 8'h67;
		16'h637B: out_word = 8'h23;
		16'h637C: out_word = 8'h1C;
		16'h637D: out_word = 8'hED;
		16'h637E: out_word = 8'h53;
		16'h637F: out_word = 8'hD7;
		16'h6380: out_word = 8'h5C;
		16'h6381: out_word = 8'hCD;
		16'h6382: out_word = 8'h9A;
		16'h6383: out_word = 8'h22;
		16'h6384: out_word = 8'hCD;
		16'h6385: out_word = 8'h70;
		16'h6386: out_word = 8'h29;
		16'h6387: out_word = 8'h0E;
		16'h6388: out_word = 8'h10;
		16'h6389: out_word = 8'hEF;
		16'h638A: out_word = 8'hEB;
		16'h638B: out_word = 8'h21;
		16'h638C: out_word = 8'hDD;
		16'h638D: out_word = 8'h5C;
		16'h638E: out_word = 8'h01;
		16'h638F: out_word = 8'h10;
		16'h6390: out_word = 8'h00;
		16'h6391: out_word = 8'hED;
		16'h6392: out_word = 8'hB0;
		16'h6393: out_word = 8'h0E;
		16'h6394: out_word = 8'h0C;
		16'h6395: out_word = 8'hEF;
		16'h6396: out_word = 8'h3A;
		16'h6397: out_word = 8'h1E;
		16'h6398: out_word = 8'h5D;
		16'h6399: out_word = 8'h77;
		16'h639A: out_word = 8'hC9;
		16'h639B: out_word = 8'h0E;
		16'h639C: out_word = 8'h0D;
		16'h639D: out_word = 8'hEF;
		16'h639E: out_word = 8'h34;
		16'h639F: out_word = 8'hC0;
		16'h63A0: out_word = 8'h23;
		16'h63A1: out_word = 8'h34;
		16'h63A2: out_word = 8'hE5;
		16'h63A3: out_word = 8'hCD;
		16'h63A4: out_word = 8'h43;
		16'h63A5: out_word = 8'h24;
		16'h63A6: out_word = 8'h0E;
		16'h63A7: out_word = 8'h23;
		16'h63A8: out_word = 8'hEF;
		16'h63A9: out_word = 8'h7E;
		16'h63AA: out_word = 8'hB7;
		16'h63AB: out_word = 8'h28;
		16'h63AC: out_word = 8'h09;
		16'h63AD: out_word = 8'hE1;
		16'h63AE: out_word = 8'hE5;
		16'h63AF: out_word = 8'h35;
		16'h63B0: out_word = 8'hCD;
		16'h63B1: out_word = 8'hFC;
		16'h63B2: out_word = 8'h23;
		16'h63B3: out_word = 8'hE1;
		16'h63B4: out_word = 8'hE5;
		16'h63B5: out_word = 8'h34;
		16'h63B6: out_word = 8'hCD;
		16'h63B7: out_word = 8'h18;
		16'h63B8: out_word = 8'h24;
		16'h63B9: out_word = 8'hE1;
		16'h63BA: out_word = 8'h3E;
		16'h63BB: out_word = 8'h10;
		16'h63BC: out_word = 8'hBE;
		16'h63BD: out_word = 8'hCC;
		16'h63BE: out_word = 8'hC1;
		16'h63BF: out_word = 8'h23;
		16'h63C0: out_word = 8'hC9;
		16'h63C1: out_word = 8'hCD;
		16'h63C2: out_word = 8'hCF;
		16'h63C3: out_word = 8'h23;
		16'h63C4: out_word = 8'hF5;
		16'h63C5: out_word = 8'hCD;
		16'h63C6: out_word = 8'h70;
		16'h63C7: out_word = 8'h29;
		16'h63C8: out_word = 8'hF1;
		16'h63C9: out_word = 8'hC2;
		16'h63CA: out_word = 8'h92;
		16'h63CB: out_word = 8'h24;
		16'h63CC: out_word = 8'hC3;
		16'h63CD: out_word = 8'h18;
		16'h63CE: out_word = 8'h24;
		16'h63CF: out_word = 8'h36;
		16'h63D0: out_word = 8'h00;
		16'h63D1: out_word = 8'h0E;
		16'h63D2: out_word = 8'h19;
		16'h63D3: out_word = 8'hEF;
		16'h63D4: out_word = 8'h34;
		16'h63D5: out_word = 8'h0E;
		16'h63D6: out_word = 8'h10;
		16'h63D7: out_word = 8'hEF;
		16'h63D8: out_word = 8'h11;
		16'h63D9: out_word = 8'hDD;
		16'h63DA: out_word = 8'h5C;
		16'h63DB: out_word = 8'h01;
		16'h63DC: out_word = 8'h10;
		16'h63DD: out_word = 8'h00;
		16'h63DE: out_word = 8'hED;
		16'h63DF: out_word = 8'hB0;
		16'h63E0: out_word = 8'hCD;
		16'h63E1: out_word = 8'hB3;
		16'h63E2: out_word = 8'h1C;
		16'h63E3: out_word = 8'hC0;
		16'h63E4: out_word = 8'hCD;
		16'h63E5: out_word = 8'h5D;
		16'h63E6: out_word = 8'h16;
		16'h63E7: out_word = 8'h0E;
		16'h63E8: out_word = 8'h10;
		16'h63E9: out_word = 8'hEF;
		16'h63EA: out_word = 8'hEB;
		16'h63EB: out_word = 8'h21;
		16'h63EC: out_word = 8'hDD;
		16'h63ED: out_word = 8'h5C;
		16'h63EE: out_word = 8'h01;
		16'h63EF: out_word = 8'h10;
		16'h63F0: out_word = 8'h00;
		16'h63F1: out_word = 8'hED;
		16'h63F2: out_word = 8'hB0;
		16'h63F3: out_word = 8'h0E;
		16'h63F4: out_word = 8'h0C;
		16'h63F5: out_word = 8'hEF;
		16'h63F6: out_word = 8'h3A;
		16'h63F7: out_word = 8'h1E;
		16'h63F8: out_word = 8'h5D;
		16'h63F9: out_word = 8'h77;
		16'h63FA: out_word = 8'hAF;
		16'h63FB: out_word = 8'hC9;
		16'h63FC: out_word = 8'hCD;
		16'h63FD: out_word = 8'h23;
		16'h63FE: out_word = 8'h24;
		16'h63FF: out_word = 8'hCD;
		16'h6400: out_word = 8'h21;
		16'h6401: out_word = 8'h23;
		16'h6402: out_word = 8'h06;
		16'h6403: out_word = 8'h01;
		16'h6404: out_word = 8'hCD;
		16'h6405: out_word = 8'h4D;
		16'h6406: out_word = 8'h1E;
		16'h6407: out_word = 8'h0E;
		16'h6408: out_word = 8'h0F;
		16'h6409: out_word = 8'hEF;
		16'h640A: out_word = 8'h7E;
		16'h640B: out_word = 8'hFE;
		16'h640C: out_word = 8'h7F;
		16'h640D: out_word = 8'hC8;
		16'h640E: out_word = 8'hCD;
		16'h640F: out_word = 8'h21;
		16'h6410: out_word = 8'h23;
		16'h6411: out_word = 8'hAF;
		16'h6412: out_word = 8'h47;
		16'h6413: out_word = 8'h77;
		16'h6414: out_word = 8'h23;
		16'h6415: out_word = 8'h10;
		16'h6416: out_word = 8'hFC;
		16'h6417: out_word = 8'hC9;
		16'h6418: out_word = 8'hCD;
		16'h6419: out_word = 8'h23;
		16'h641A: out_word = 8'h24;
		16'h641B: out_word = 8'hCD;
		16'h641C: out_word = 8'h21;
		16'h641D: out_word = 8'h23;
		16'h641E: out_word = 8'h06;
		16'h641F: out_word = 8'h01;
		16'h6420: out_word = 8'hC3;
		16'h6421: out_word = 8'h3D;
		16'h6422: out_word = 8'h1E;
		16'h6423: out_word = 8'h2A;
		16'h6424: out_word = 8'h51;
		16'h6425: out_word = 8'h5C;
		16'h6426: out_word = 8'h01;
		16'h6427: out_word = 8'h1E;
		16'h6428: out_word = 8'h00;
		16'h6429: out_word = 8'h09;
		16'h642A: out_word = 8'h5E;
		16'h642B: out_word = 8'h23;
		16'h642C: out_word = 8'h56;
		16'h642D: out_word = 8'h0E;
		16'h642E: out_word = 8'h0E;
		16'h642F: out_word = 8'hEF;
		16'h6430: out_word = 8'h46;
		16'h6431: out_word = 8'h05;
		16'h6432: out_word = 8'h04;
		16'h6433: out_word = 8'hF5;
		16'h6434: out_word = 8'h3E;
		16'h6435: out_word = 8'h10;
		16'h6436: out_word = 8'h28;
		16'h6437: out_word = 8'h09;
		16'h6438: out_word = 8'h1C;
		16'h6439: out_word = 8'hBB;
		16'h643A: out_word = 8'h20;
		16'h643B: out_word = 8'h03;
		16'h643C: out_word = 8'h1E;
		16'h643D: out_word = 8'h00;
		16'h643E: out_word = 8'h14;
		16'h643F: out_word = 8'h10;
		16'h6440: out_word = 8'hF7;
		16'h6441: out_word = 8'hF1;
		16'h6442: out_word = 8'hC9;
		16'h6443: out_word = 8'h0E;
		16'h6444: out_word = 8'h0B;
		16'h6445: out_word = 8'hEF;
		16'h6446: out_word = 8'h7E;
		16'h6447: out_word = 8'hC3;
		16'h6448: out_word = 8'hCB;
		16'h6449: out_word = 8'h3D;
		16'h644A: out_word = 8'h21;
		16'h644B: out_word = 8'hC2;
		16'h644C: out_word = 8'h5C;
		16'h644D: out_word = 8'hE5;
		16'h644E: out_word = 8'h21;
		16'h644F: out_word = 8'hF1;
		16'h6450: out_word = 8'h20;
		16'h6451: out_word = 8'hE5;
		16'h6452: out_word = 8'hF5;
		16'h6453: out_word = 8'hCD;
		16'h6454: out_word = 8'hF1;
		16'h6455: out_word = 8'h20;
		16'h6456: out_word = 8'h3E;
		16'h6457: out_word = 8'h0A;
		16'h6458: out_word = 8'h32;
		16'h6459: out_word = 8'h06;
		16'h645A: out_word = 8'h5D;
		16'h645B: out_word = 8'hF1;
		16'h645C: out_word = 8'hCD;
		16'h645D: out_word = 8'hA2;
		16'h645E: out_word = 8'h24;
		16'h645F: out_word = 8'hF5;
		16'h6460: out_word = 8'hCD;
		16'h6461: out_word = 8'h50;
		16'h6462: out_word = 8'h26;
		16'h6463: out_word = 8'hCA;
		16'h6464: out_word = 8'h9E;
		16'h6465: out_word = 8'h24;
		16'h6466: out_word = 8'hF1;
		16'h6467: out_word = 8'hCD;
		16'h6468: out_word = 8'h17;
		16'h6469: out_word = 8'h23;
		16'h646A: out_word = 8'h77;
		16'h646B: out_word = 8'hC3;
		16'h646C: out_word = 8'h2A;
		16'h646D: out_word = 8'h23;
		16'h646E: out_word = 8'h0E;
		16'h646F: out_word = 8'h0D;
		16'h6470: out_word = 8'hEF;
		16'h6471: out_word = 8'h7E;
		16'h6472: out_word = 8'h01;
		16'h6473: out_word = 8'h0E;
		16'h6474: out_word = 8'h00;
		16'h6475: out_word = 8'h09;
		16'h6476: out_word = 8'hBE;
		16'h6477: out_word = 8'hC0;
		16'h6478: out_word = 8'h0E;
		16'h6479: out_word = 8'h0E;
		16'h647A: out_word = 8'hEF;
		16'h647B: out_word = 8'h7E;
		16'h647C: out_word = 8'h01;
		16'h647D: out_word = 8'h0E;
		16'h647E: out_word = 8'h00;
		16'h647F: out_word = 8'h09;
		16'h6480: out_word = 8'hBE;
		16'h6481: out_word = 8'hC0;
		16'h6482: out_word = 8'h21;
		16'h6483: out_word = 8'hB6;
		16'h6484: out_word = 8'h5C;
		16'h6485: out_word = 8'h7E;
		16'h6486: out_word = 8'hFE;
		16'h6487: out_word = 8'hF4;
		16'h6488: out_word = 8'h28;
		16'h6489: out_word = 8'h08;
		16'h648A: out_word = 8'hCB;
		16'h648B: out_word = 8'h66;
		16'h648C: out_word = 8'h28;
		16'h648D: out_word = 8'h04;
		16'h648E: out_word = 8'hF6;
		16'h648F: out_word = 8'h01;
		16'h6490: out_word = 8'hE1;
		16'h6491: out_word = 8'hC9;
		16'h6492: out_word = 8'h3E;
		16'h6493: out_word = 8'h07;
		16'h6494: out_word = 8'h32;
		16'h6495: out_word = 8'h3A;
		16'h6496: out_word = 8'h5C;
		16'h6497: out_word = 8'hCD;
		16'h6498: out_word = 8'hE5;
		16'h6499: out_word = 8'h20;
		16'h649A: out_word = 8'hE7;
		16'h649B: out_word = 8'h58;
		16'h649C: out_word = 8'h00;
		16'h649D: out_word = 8'hC9;
		16'h649E: out_word = 8'h3E;
		16'h649F: out_word = 8'h17;
		16'h64A0: out_word = 8'h18;
		16'h64A1: out_word = 8'hF2;
		16'h64A2: out_word = 8'h57;
		16'h64A3: out_word = 8'h0E;
		16'h64A4: out_word = 8'h0F;
		16'h64A5: out_word = 8'hEF;
		16'h64A6: out_word = 8'h7E;
		16'h64A7: out_word = 8'hFE;
		16'h64A8: out_word = 8'h7F;
		16'h64A9: out_word = 8'h7A;
		16'h64AA: out_word = 8'hC0;
		16'h64AB: out_word = 8'h01;
		16'h64AC: out_word = 8'h13;
		16'h64AD: out_word = 8'h00;
		16'h64AE: out_word = 8'h09;
		16'h64AF: out_word = 8'h7E;
		16'h64B0: out_word = 8'hB7;
		16'h64B1: out_word = 8'h7A;
		16'h64B2: out_word = 8'h20;
		16'h64B3: out_word = 8'h21;
		16'h64B4: out_word = 8'h2B;
		16'h64B5: out_word = 8'h7E;
		16'h64B6: out_word = 8'hB7;
		16'h64B7: out_word = 8'h20;
		16'h64B8: out_word = 8'h09;
		16'h64B9: out_word = 8'hC5;
		16'h64BA: out_word = 8'hE5;
		16'h64BB: out_word = 8'hD5;
		16'h64BC: out_word = 8'hCD;
		16'h64BD: out_word = 8'hF8;
		16'h64BE: out_word = 8'h24;
		16'h64BF: out_word = 8'hD1;
		16'h64C0: out_word = 8'hE1;
		16'h64C1: out_word = 8'hC1;
		16'h64C2: out_word = 8'h4E;
		16'h64C3: out_word = 8'h7A;
		16'h64C4: out_word = 8'hEB;
		16'h64C5: out_word = 8'h2A;
		16'h64C6: out_word = 8'hCF;
		16'h64C7: out_word = 8'h5C;
		16'h64C8: out_word = 8'h09;
		16'h64C9: out_word = 8'hFE;
		16'h64CA: out_word = 8'h06;
		16'h64CB: out_word = 8'h77;
		16'h64CC: out_word = 8'hCC;
		16'h64CD: out_word = 8'h04;
		16'h64CE: out_word = 8'h25;
		16'h64CF: out_word = 8'h0E;
		16'h64D0: out_word = 8'h21;
		16'h64D1: out_word = 8'hEF;
		16'h64D2: out_word = 8'h34;
		16'h64D3: out_word = 8'hE1;
		16'h64D4: out_word = 8'hC9;
		16'h64D5: out_word = 8'h2B;
		16'h64D6: out_word = 8'h7E;
		16'h64D7: out_word = 8'h2B;
		16'h64D8: out_word = 8'h3C;
		16'h64D9: out_word = 8'hBE;
		16'h64DA: out_word = 8'h23;
		16'h64DB: out_word = 8'h34;
		16'h64DC: out_word = 8'hE5;
		16'h64DD: out_word = 8'hF5;
		16'h64DE: out_word = 8'h0E;
		16'h64DF: out_word = 8'h23;
		16'h64E0: out_word = 8'hEF;
		16'h64E1: out_word = 8'h36;
		16'h64E2: out_word = 8'hFF;
		16'h64E3: out_word = 8'hF1;
		16'h64E4: out_word = 8'hE1;
		16'h64E5: out_word = 8'h38;
		16'h64E6: out_word = 8'h07;
		16'h64E7: out_word = 8'h7A;
		16'h64E8: out_word = 8'hFE;
		16'h64E9: out_word = 8'h0D;
		16'h64EA: out_word = 8'h28;
		16'h64EB: out_word = 8'h06;
		16'h64EC: out_word = 8'hC1;
		16'h64ED: out_word = 8'hC9;
		16'h64EE: out_word = 8'h7A;
		16'h64EF: out_word = 8'hFE;
		16'h64F0: out_word = 8'h0D;
		16'h64F1: out_word = 8'hC0;
		16'h64F2: out_word = 8'hAF;
		16'h64F3: out_word = 8'h77;
		16'h64F4: out_word = 8'h23;
		16'h64F5: out_word = 8'h77;
		16'h64F6: out_word = 8'h7A;
		16'h64F7: out_word = 8'hC9;
		16'h64F8: out_word = 8'h2A;
		16'h64F9: out_word = 8'h61;
		16'h64FA: out_word = 8'h5C;
		16'h64FB: out_word = 8'h22;
		16'h64FC: out_word = 8'hCF;
		16'h64FD: out_word = 8'h5C;
		16'h64FE: out_word = 8'h01;
		16'h64FF: out_word = 8'h10;
		16'h6500: out_word = 8'h00;
		16'h6501: out_word = 8'hC3;
		16'h6502: out_word = 8'h23;
		16'h6503: out_word = 8'h1E;
		16'h6504: out_word = 8'h36;
		16'h6505: out_word = 8'h0D;
		16'h6506: out_word = 8'h2A;
		16'h6507: out_word = 8'h5D;
		16'h6508: out_word = 8'h5C;
		16'h6509: out_word = 8'h22;
		16'h650A: out_word = 8'hD7;
		16'h650B: out_word = 8'h5C;
		16'h650C: out_word = 8'h2A;
		16'h650D: out_word = 8'hCF;
		16'h650E: out_word = 8'h5C;
		16'h650F: out_word = 8'h22;
		16'h6510: out_word = 8'h5D;
		16'h6511: out_word = 8'h5C;
		16'h6512: out_word = 8'h21;
		16'h6513: out_word = 8'h3B;
		16'h6514: out_word = 8'h5C;
		16'h6515: out_word = 8'hCB;
		16'h6516: out_word = 8'hBE;
		16'h6517: out_word = 8'hCD;
		16'h6518: out_word = 8'hC1;
		16'h6519: out_word = 8'h1D;
		16'h651A: out_word = 8'h21;
		16'h651B: out_word = 8'h3B;
		16'h651C: out_word = 8'h5C;
		16'h651D: out_word = 8'hCB;
		16'h651E: out_word = 8'hFE;
		16'h651F: out_word = 8'h2A;
		16'h6520: out_word = 8'hCF;
		16'h6521: out_word = 8'h5C;
		16'h6522: out_word = 8'h22;
		16'h6523: out_word = 8'h5D;
		16'h6524: out_word = 8'h5C;
		16'h6525: out_word = 8'hCD;
		16'h6526: out_word = 8'hC1;
		16'h6527: out_word = 8'h1D;
		16'h6528: out_word = 8'hCD;
		16'h6529: out_word = 8'hB9;
		16'h652A: out_word = 8'h1D;
		16'h652B: out_word = 8'hC5;
		16'h652C: out_word = 8'hD1;
		16'h652D: out_word = 8'h0E;
		16'h652E: out_word = 8'h20;
		16'h652F: out_word = 8'hEF;
		16'h6530: out_word = 8'h46;
		16'h6531: out_word = 8'hAF;
		16'h6532: out_word = 8'h21;
		16'h6533: out_word = 8'h00;
		16'h6534: out_word = 8'h00;
		16'h6535: out_word = 8'h22;
		16'h6536: out_word = 8'hDB;
		16'h6537: out_word = 8'h5C;
		16'h6538: out_word = 8'h19;
		16'h6539: out_word = 8'h30;
		16'h653A: out_word = 8'h09;
		16'h653B: out_word = 8'hE5;
		16'h653C: out_word = 8'h2A;
		16'h653D: out_word = 8'hDB;
		16'h653E: out_word = 8'h5C;
		16'h653F: out_word = 8'h23;
		16'h6540: out_word = 8'h22;
		16'h6541: out_word = 8'hDB;
		16'h6542: out_word = 8'h5C;
		16'h6543: out_word = 8'hE1;
		16'h6544: out_word = 8'h10;
		16'h6545: out_word = 8'hF2;
		16'h6546: out_word = 8'h22;
		16'h6547: out_word = 8'hD9;
		16'h6548: out_word = 8'h5C;
		16'h6549: out_word = 8'h3A;
		16'h654A: out_word = 8'hDB;
		16'h654B: out_word = 8'h5C;
		16'h654C: out_word = 8'h21;
		16'h654D: out_word = 8'hDA;
		16'h654E: out_word = 8'h5C;
		16'h654F: out_word = 8'hED;
		16'h6550: out_word = 8'h67;
		16'h6551: out_word = 8'hE6;
		16'h6552: out_word = 8'h0F;
		16'h6553: out_word = 8'h32;
		16'h6554: out_word = 8'hDB;
		16'h6555: out_word = 8'h5C;
		16'h6556: out_word = 8'h2A;
		16'h6557: out_word = 8'hD7;
		16'h6558: out_word = 8'h5C;
		16'h6559: out_word = 8'h22;
		16'h655A: out_word = 8'h5D;
		16'h655B: out_word = 8'h5C;
		16'h655C: out_word = 8'hCD;
		16'h655D: out_word = 8'h68;
		16'h655E: out_word = 8'h25;
		16'h655F: out_word = 8'h0E;
		16'h6560: out_word = 8'h21;
		16'h6561: out_word = 8'hEF;
		16'h6562: out_word = 8'h3E;
		16'h6563: out_word = 8'hFF;
		16'h6564: out_word = 8'h77;
		16'h6565: out_word = 8'h23;
		16'h6566: out_word = 8'h77;
		16'h6567: out_word = 8'hC9;
		16'h6568: out_word = 8'h0E;
		16'h6569: out_word = 8'h19;
		16'h656A: out_word = 8'hEF;
		16'h656B: out_word = 8'h3A;
		16'h656C: out_word = 8'hDA;
		16'h656D: out_word = 8'h5C;
		16'h656E: out_word = 8'hBE;
		16'h656F: out_word = 8'hC2;
		16'h6570: out_word = 8'h84;
		16'h6571: out_word = 8'h25;
		16'h6572: out_word = 8'h0E;
		16'h6573: out_word = 8'h0E;
		16'h6574: out_word = 8'hEF;
		16'h6575: out_word = 8'h3A;
		16'h6576: out_word = 8'hDB;
		16'h6577: out_word = 8'h5C;
		16'h6578: out_word = 8'hBE;
		16'h6579: out_word = 8'hC2;
		16'h657A: out_word = 8'hA7;
		16'h657B: out_word = 8'h25;
		16'h657C: out_word = 8'h0E;
		16'h657D: out_word = 8'h0D;
		16'h657E: out_word = 8'hEF;
		16'h657F: out_word = 8'h3A;
		16'h6580: out_word = 8'hD9;
		16'h6581: out_word = 8'h5C;
		16'h6582: out_word = 8'h77;
		16'h6583: out_word = 8'hC9;
		16'h6584: out_word = 8'hCD;
		16'h6585: out_word = 8'hCA;
		16'h6586: out_word = 8'h25;
		16'h6587: out_word = 8'hC4;
		16'h6588: out_word = 8'hC3;
		16'h6589: out_word = 8'h25;
		16'h658A: out_word = 8'h3A;
		16'h658B: out_word = 8'hDA;
		16'h658C: out_word = 8'h5C;
		16'h658D: out_word = 8'h0E;
		16'h658E: out_word = 8'h19;
		16'h658F: out_word = 8'hEF;
		16'h6590: out_word = 8'h77;
		16'h6591: out_word = 8'h0E;
		16'h6592: out_word = 8'h10;
		16'h6593: out_word = 8'hEF;
		16'h6594: out_word = 8'h11;
		16'h6595: out_word = 8'hDD;
		16'h6596: out_word = 8'h5C;
		16'h6597: out_word = 8'h01;
		16'h6598: out_word = 8'h10;
		16'h6599: out_word = 8'h00;
		16'h659A: out_word = 8'hED;
		16'h659B: out_word = 8'hB0;
		16'h659C: out_word = 8'hCD;
		16'h659D: out_word = 8'hB3;
		16'h659E: out_word = 8'h1C;
		16'h659F: out_word = 8'hC2;
		16'h65A0: out_word = 8'hD2;
		16'h65A1: out_word = 8'h25;
		16'h65A2: out_word = 8'hCD;
		16'h65A3: out_word = 8'hE4;
		16'h65A4: out_word = 8'h23;
		16'h65A5: out_word = 8'h18;
		16'h65A6: out_word = 8'h06;
		16'h65A7: out_word = 8'hCD;
		16'h65A8: out_word = 8'hCA;
		16'h65A9: out_word = 8'h25;
		16'h65AA: out_word = 8'hC4;
		16'h65AB: out_word = 8'hC3;
		16'h65AC: out_word = 8'h25;
		16'h65AD: out_word = 8'h3A;
		16'h65AE: out_word = 8'hDB;
		16'h65AF: out_word = 8'h5C;
		16'h65B0: out_word = 8'h0E;
		16'h65B1: out_word = 8'h0E;
		16'h65B2: out_word = 8'hEF;
		16'h65B3: out_word = 8'h77;
		16'h65B4: out_word = 8'hE5;
		16'h65B5: out_word = 8'hCD;
		16'h65B6: out_word = 8'h43;
		16'h65B7: out_word = 8'h24;
		16'h65B8: out_word = 8'hCD;
		16'h65B9: out_word = 8'h18;
		16'h65BA: out_word = 8'h24;
		16'h65BB: out_word = 8'hE1;
		16'h65BC: out_word = 8'h2B;
		16'h65BD: out_word = 8'h3A;
		16'h65BE: out_word = 8'hD9;
		16'h65BF: out_word = 8'h5C;
		16'h65C0: out_word = 8'h77;
		16'h65C1: out_word = 8'h18;
		16'h65C2: out_word = 8'hB9;
		16'h65C3: out_word = 8'hCD;
		16'h65C4: out_word = 8'h43;
		16'h65C5: out_word = 8'h24;
		16'h65C6: out_word = 8'hCD;
		16'h65C7: out_word = 8'hFC;
		16'h65C8: out_word = 8'h23;
		16'h65C9: out_word = 8'hC9;
		16'h65CA: out_word = 8'h0E;
		16'h65CB: out_word = 8'h23;
		16'h65CC: out_word = 8'hEF;
		16'h65CD: out_word = 8'h7E;
		16'h65CE: out_word = 8'hB7;
		16'h65CF: out_word = 8'h36;
		16'h65D0: out_word = 8'h00;
		16'h65D1: out_word = 8'hC9;
		16'h65D2: out_word = 8'h2A;
		16'h65D3: out_word = 8'hDA;
		16'h65D4: out_word = 8'h5C;
		16'h65D5: out_word = 8'h26;
		16'h65D6: out_word = 8'h20;
		16'h65D7: out_word = 8'h22;
		16'h65D8: out_word = 8'hD7;
		16'h65D9: out_word = 8'h5C;
		16'h65DA: out_word = 8'h2A;
		16'h65DB: out_word = 8'hD9;
		16'h65DC: out_word = 8'h5C;
		16'h65DD: out_word = 8'hE5;
		16'h65DE: out_word = 8'h2A;
		16'h65DF: out_word = 8'hDB;
		16'h65E0: out_word = 8'h5C;
		16'h65E1: out_word = 8'hE5;
		16'h65E2: out_word = 8'hCD;
		16'h65E3: out_word = 8'h81;
		16'h65E4: out_word = 8'h23;
		16'h65E5: out_word = 8'hE1;
		16'h65E6: out_word = 8'h22;
		16'h65E7: out_word = 8'hDB;
		16'h65E8: out_word = 8'h5C;
		16'h65E9: out_word = 8'hE1;
		16'h65EA: out_word = 8'h22;
		16'h65EB: out_word = 8'hD9;
		16'h65EC: out_word = 8'h5C;
		16'h65ED: out_word = 8'h18;
		16'h65EE: out_word = 8'hBE;
		16'h65EF: out_word = 8'hCD;
		16'h65F0: out_word = 8'hF1;
		16'h65F1: out_word = 8'h20;
		16'h65F2: out_word = 8'h21;
		16'h65F3: out_word = 8'h3C;
		16'h65F4: out_word = 8'h5C;
		16'h65F5: out_word = 8'hCB;
		16'h65F6: out_word = 8'h9E;
		16'h65F7: out_word = 8'h2A;
		16'h65F8: out_word = 8'h3D;
		16'h65F9: out_word = 8'h5C;
		16'h65FA: out_word = 8'h5E;
		16'h65FB: out_word = 8'h23;
		16'h65FC: out_word = 8'h56;
		16'h65FD: out_word = 8'hB7;
		16'h65FE: out_word = 8'h21;
		16'h65FF: out_word = 8'h7F;
		16'h6600: out_word = 8'h10;
		16'h6601: out_word = 8'hED;
		16'h6602: out_word = 8'h52;
		16'h6603: out_word = 8'h20;
		16'h6604: out_word = 8'h21;
		16'h6605: out_word = 8'hED;
		16'h6606: out_word = 8'h7B;
		16'h6607: out_word = 8'h3D;
		16'h6608: out_word = 8'h5C;
		16'h6609: out_word = 8'hD1;
		16'h660A: out_word = 8'hD1;
		16'h660B: out_word = 8'hED;
		16'h660C: out_word = 8'h53;
		16'h660D: out_word = 8'h3D;
		16'h660E: out_word = 8'h5C;
		16'h660F: out_word = 8'hCD;
		16'h6610: out_word = 8'h2B;
		16'h6611: out_word = 8'h26;
		16'h6612: out_word = 8'h38;
		16'h6613: out_word = 8'h09;
		16'h6614: out_word = 8'h21;
		16'h6615: out_word = 8'hC2;
		16'h6616: out_word = 8'h5C;
		16'h6617: out_word = 8'hE5;
		16'h6618: out_word = 8'h21;
		16'h6619: out_word = 8'hE5;
		16'h661A: out_word = 8'h20;
		16'h661B: out_word = 8'hE5;
		16'h661C: out_word = 8'hC9;
		16'h661D: out_word = 8'hFE;
		16'h661E: out_word = 8'h0D;
		16'h661F: out_word = 8'h28;
		16'h6620: out_word = 8'hF3;
		16'h6621: out_word = 8'hE7;
		16'h6622: out_word = 8'h85;
		16'h6623: out_word = 8'h0F;
		16'h6624: out_word = 8'h18;
		16'h6625: out_word = 8'hE9;
		16'h6626: out_word = 8'hCD;
		16'h6627: out_word = 8'h2B;
		16'h6628: out_word = 8'h26;
		16'h6629: out_word = 8'h18;
		16'h662A: out_word = 8'hE9;
		16'h662B: out_word = 8'h3E;
		16'h662C: out_word = 8'h0A;
		16'h662D: out_word = 8'h32;
		16'h662E: out_word = 8'h06;
		16'h662F: out_word = 8'h5D;
		16'h6630: out_word = 8'hCD;
		16'h6631: out_word = 8'h50;
		16'h6632: out_word = 8'h26;
		16'h6633: out_word = 8'h28;
		16'h6634: out_word = 8'h0D;
		16'h6635: out_word = 8'hFE;
		16'h6636: out_word = 8'h7F;
		16'h6637: out_word = 8'hC2;
		16'h6638: out_word = 8'h9E;
		16'h6639: out_word = 8'h24;
		16'h663A: out_word = 8'h01;
		16'h663B: out_word = 8'h13;
		16'h663C: out_word = 8'h00;
		16'h663D: out_word = 8'h09;
		16'h663E: out_word = 8'h36;
		16'h663F: out_word = 8'h00;
		16'h6640: out_word = 8'h18;
		16'h6641: out_word = 8'h03;
		16'h6642: out_word = 8'hCD;
		16'h6643: out_word = 8'h6E;
		16'h6644: out_word = 8'h24;
		16'h6645: out_word = 8'hCD;
		16'h6646: out_word = 8'h17;
		16'h6647: out_word = 8'h23;
		16'h6648: out_word = 8'h7E;
		16'h6649: out_word = 8'hF5;
		16'h664A: out_word = 8'hCD;
		16'h664B: out_word = 8'h9B;
		16'h664C: out_word = 8'h23;
		16'h664D: out_word = 8'hF1;
		16'h664E: out_word = 8'h37;
		16'h664F: out_word = 8'hC9;
		16'h6650: out_word = 8'h0E;
		16'h6651: out_word = 8'h0F;
		16'h6652: out_word = 8'hEF;
		16'h6653: out_word = 8'h7E;
		16'h6654: out_word = 8'hB7;
		16'h6655: out_word = 8'hC9;
		16'h6656: out_word = 8'h2A;
		16'h6657: out_word = 8'h11;
		16'h6658: out_word = 8'h5D;
		16'h6659: out_word = 8'h22;
		16'h665A: out_word = 8'h5D;
		16'h665B: out_word = 8'h5C;
		16'h665C: out_word = 8'hCD;
		16'h665D: out_word = 8'h0B;
		16'h665E: out_word = 8'h1E;
		16'h665F: out_word = 8'hCD;
		16'h6660: out_word = 8'h75;
		16'h6661: out_word = 8'h1D;
		16'h6662: out_word = 8'h3A;
		16'h6663: out_word = 8'hDB;
		16'h6664: out_word = 8'h5C;
		16'h6665: out_word = 8'hE7;
		16'h6666: out_word = 8'h27;
		16'h6667: out_word = 8'h17;
		16'h6668: out_word = 8'h78;
		16'h6669: out_word = 8'hB1;
		16'h666A: out_word = 8'hCA;
		16'h666B: out_word = 8'hD3;
		16'h666C: out_word = 8'h01;
		16'h666D: out_word = 8'hE5;
		16'h666E: out_word = 8'h2A;
		16'h666F: out_word = 8'h4F;
		16'h6670: out_word = 8'h5C;
		16'h6671: out_word = 8'h09;
		16'h6672: out_word = 8'h7E;
		16'h6673: out_word = 8'h21;
		16'h6674: out_word = 8'h0E;
		16'h6675: out_word = 8'h3D;
		16'h6676: out_word = 8'hBC;
		16'h6677: out_word = 8'hE1;
		16'h6678: out_word = 8'hC2;
		16'h6679: out_word = 8'h28;
		16'h667A: out_word = 8'h22;
		16'h667B: out_word = 8'h36;
		16'h667C: out_word = 8'h00;
		16'h667D: out_word = 8'h23;
		16'h667E: out_word = 8'h36;
		16'h667F: out_word = 8'h00;
		16'h6680: out_word = 8'hED;
		16'h6681: out_word = 8'h43;
		16'h6682: out_word = 8'hD9;
		16'h6683: out_word = 8'h5C;
		16'h6684: out_word = 8'h2A;
		16'h6685: out_word = 8'h4F;
		16'h6686: out_word = 8'h5C;
		16'h6687: out_word = 8'h09;
		16'h6688: out_word = 8'h2B;
		16'h6689: out_word = 8'h22;
		16'h668A: out_word = 8'hD7;
		16'h668B: out_word = 8'h5C;
		16'h668C: out_word = 8'hCD;
		16'h668D: out_word = 8'hCE;
		16'h668E: out_word = 8'h26;
		16'h668F: out_word = 8'h2A;
		16'h6690: out_word = 8'hD7;
		16'h6691: out_word = 8'h5C;
		16'h6692: out_word = 8'h01;
		16'h6693: out_word = 8'h24;
		16'h6694: out_word = 8'h01;
		16'h6695: out_word = 8'hCD;
		16'h6696: out_word = 8'h2E;
		16'h6697: out_word = 8'h1E;
		16'h6698: out_word = 8'h21;
		16'h6699: out_word = 8'h10;
		16'h669A: out_word = 8'h5C;
		16'h669B: out_word = 8'h06;
		16'h669C: out_word = 8'h10;
		16'h669D: out_word = 8'hC5;
		16'h669E: out_word = 8'hED;
		16'h669F: out_word = 8'h4B;
		16'h66A0: out_word = 8'hD9;
		16'h66A1: out_word = 8'h5C;
		16'h66A2: out_word = 8'h5E;
		16'h66A3: out_word = 8'h23;
		16'h66A4: out_word = 8'h56;
		16'h66A5: out_word = 8'hEB;
		16'h66A6: out_word = 8'hED;
		16'h66A7: out_word = 8'h42;
		16'h66A8: out_word = 8'hEB;
		16'h66A9: out_word = 8'h38;
		16'h66AA: out_word = 8'h11;
		16'h66AB: out_word = 8'h56;
		16'h66AC: out_word = 8'h2B;
		16'h66AD: out_word = 8'h5E;
		16'h66AE: out_word = 8'h23;
		16'h66AF: out_word = 8'hE5;
		16'h66B0: out_word = 8'hEB;
		16'h66B1: out_word = 8'h01;
		16'h66B2: out_word = 8'h24;
		16'h66B3: out_word = 8'h01;
		16'h66B4: out_word = 8'hED;
		16'h66B5: out_word = 8'h42;
		16'h66B6: out_word = 8'hEB;
		16'h66B7: out_word = 8'hE1;
		16'h66B8: out_word = 8'h72;
		16'h66B9: out_word = 8'h2B;
		16'h66BA: out_word = 8'h73;
		16'h66BB: out_word = 8'h23;
		16'h66BC: out_word = 8'h23;
		16'h66BD: out_word = 8'hC1;
		16'h66BE: out_word = 8'h10;
		16'h66BF: out_word = 8'hDD;
		16'h66C0: out_word = 8'h2A;
		16'h66C1: out_word = 8'h11;
		16'h66C2: out_word = 8'h5D;
		16'h66C3: out_word = 8'h01;
		16'h66C4: out_word = 8'h24;
		16'h66C5: out_word = 8'h01;
		16'h66C6: out_word = 8'hED;
		16'h66C7: out_word = 8'h42;
		16'h66C8: out_word = 8'h22;
		16'h66C9: out_word = 8'h11;
		16'h66CA: out_word = 8'h5D;
		16'h66CB: out_word = 8'hC3;
		16'h66CC: out_word = 8'hD3;
		16'h66CD: out_word = 8'h01;
		16'h66CE: out_word = 8'h01;
		16'h66CF: out_word = 8'h0F;
		16'h66D0: out_word = 8'h00;
		16'h66D1: out_word = 8'h09;
		16'h66D2: out_word = 8'h7E;
		16'h66D3: out_word = 8'hB7;
		16'h66D4: out_word = 8'hC8;
		16'h66D5: out_word = 8'h2A;
		16'h66D6: out_word = 8'hD7;
		16'h66D7: out_word = 8'h5C;
		16'h66D8: out_word = 8'h22;
		16'h66D9: out_word = 8'h51;
		16'h66DA: out_word = 8'h5C;
		16'h66DB: out_word = 8'hCD;
		16'h66DC: out_word = 8'hE1;
		16'h66DD: out_word = 8'h26;
		16'h66DE: out_word = 8'hC3;
		16'h66DF: out_word = 8'hFC;
		16'h66E0: out_word = 8'h23;
		16'h66E1: out_word = 8'h01;
		16'h66E2: out_word = 8'h0D;
		16'h66E3: out_word = 8'h00;
		16'h66E4: out_word = 8'h09;
		16'h66E5: out_word = 8'h5E;
		16'h66E6: out_word = 8'h23;
		16'h66E7: out_word = 8'h56;
		16'h66E8: out_word = 8'h01;
		16'h66E9: out_word = 8'h0D;
		16'h66EA: out_word = 8'h00;
		16'h66EB: out_word = 8'h09;
		16'h66EC: out_word = 8'h73;
		16'h66ED: out_word = 8'h23;
		16'h66EE: out_word = 8'h72;
		16'h66EF: out_word = 8'h0E;
		16'h66F0: out_word = 8'h10;
		16'h66F1: out_word = 8'hEF;
		16'h66F2: out_word = 8'h11;
		16'h66F3: out_word = 8'hDD;
		16'h66F4: out_word = 8'h5C;
		16'h66F5: out_word = 8'h01;
		16'h66F6: out_word = 8'h10;
		16'h66F7: out_word = 8'h00;
		16'h66F8: out_word = 8'hED;
		16'h66F9: out_word = 8'hB0;
		16'h66FA: out_word = 8'hCD;
		16'h66FB: out_word = 8'h43;
		16'h66FC: out_word = 8'h24;
		16'h66FD: out_word = 8'h0E;
		16'h66FE: out_word = 8'h0C;
		16'h66FF: out_word = 8'hEF;
		16'h6700: out_word = 8'h4E;
		16'h6701: out_word = 8'hCD;
		16'h6702: out_word = 8'h6B;
		16'h6703: out_word = 8'h16;
		16'h6704: out_word = 8'hC3;
		16'h6705: out_word = 8'h43;
		16'h6706: out_word = 8'h1E;
		16'h6707: out_word = 8'h7E;
		16'h6708: out_word = 8'hB7;
		16'h6709: out_word = 8'hC8;
		16'h670A: out_word = 8'hE6;
		16'h670B: out_word = 8'h7F;
		16'h670C: out_word = 8'hD7;
		16'h670D: out_word = 8'hCB;
		16'h670E: out_word = 8'h7E;
		16'h670F: out_word = 8'hC0;
		16'h6710: out_word = 8'h23;
		16'h6711: out_word = 8'h18;
		16'h6712: out_word = 8'hF4;
		16'h6713: out_word = 8'h1A;
		16'h6714: out_word = 8'hBE;
		16'h6715: out_word = 8'hC0;
		16'h6716: out_word = 8'h13;
		16'h6717: out_word = 8'h23;
		16'h6718: out_word = 8'h10;
		16'h6719: out_word = 8'hF9;
		16'h671A: out_word = 8'hC9;
		16'h671B: out_word = 8'h21;
		16'h671C: out_word = 8'hFC;
		16'h671D: out_word = 8'h27;
		16'h671E: out_word = 8'h3E;
		16'h671F: out_word = 8'h06;
		16'h6720: out_word = 8'hC3;
		16'h6721: out_word = 8'h4A;
		16'h6722: out_word = 8'h1C;
		16'h6723: out_word = 8'h21;
		16'h6724: out_word = 8'hED;
		16'h6725: out_word = 8'h27;
		16'h6726: out_word = 8'h3E;
		16'h6727: out_word = 8'h04;
		16'h6728: out_word = 8'hC3;
		16'h6729: out_word = 8'h4A;
		16'h672A: out_word = 8'h1C;
		16'h672B: out_word = 8'h3E;
		16'h672C: out_word = 8'h1A;
		16'h672D: out_word = 8'h18;
		16'h672E: out_word = 8'h02;
		16'h672F: out_word = 8'h3E;
		16'h6730: out_word = 8'h12;
		16'h6731: out_word = 8'h32;
		16'h6732: out_word = 8'h3A;
		16'h6733: out_word = 8'h5C;
		16'h6734: out_word = 8'hC9;
		16'h6735: out_word = 8'h3E;
		16'h6736: out_word = 8'h03;
		16'h6737: out_word = 8'h18;
		16'h6738: out_word = 8'hF8;
		16'h6739: out_word = 8'hAF;
		16'h673A: out_word = 8'h32;
		16'h673B: out_word = 8'hD8;
		16'h673C: out_word = 8'h5C;
		16'h673D: out_word = 8'h32;
		16'h673E: out_word = 8'hD6;
		16'h673F: out_word = 8'h5C;
		16'h6740: out_word = 8'hDB;
		16'h6741: out_word = 8'h1F;
		16'h6742: out_word = 8'h32;
		16'h6743: out_word = 8'hCD;
		16'h6744: out_word = 8'h5C;
		16'h6745: out_word = 8'h5A;
		16'h6746: out_word = 8'hD5;
		16'h6747: out_word = 8'h7B;
		16'h6748: out_word = 8'hD3;
		16'h6749: out_word = 8'h7F;
		16'h674A: out_word = 8'h3E;
		16'h674B: out_word = 8'h18;
		16'h674C: out_word = 8'hCD;
		16'h674D: out_word = 8'h9A;
		16'h674E: out_word = 8'h3D;
		16'h674F: out_word = 8'h3A;
		16'h6750: out_word = 8'hCD;
		16'h6751: out_word = 8'h5C;
		16'h6752: out_word = 8'hE6;
		16'h6753: out_word = 8'h80;
		16'h6754: out_word = 8'hC4;
		16'h6755: out_word = 8'hA0;
		16'h6756: out_word = 8'h3E;
		16'h6757: out_word = 8'hD1;
		16'h6758: out_word = 8'hCD;
		16'h6759: out_word = 8'h7D;
		16'h675A: out_word = 8'h20;
		16'h675B: out_word = 8'h3A;
		16'h675C: out_word = 8'hD6;
		16'h675D: out_word = 8'h5C;
		16'h675E: out_word = 8'hB7;
		16'h675F: out_word = 8'hC8;
		16'h6760: out_word = 8'h3E;
		16'h6761: out_word = 8'h07;
		16'h6762: out_word = 8'h32;
		16'h6763: out_word = 8'h0F;
		16'h6764: out_word = 8'h5D;
		16'h6765: out_word = 8'hC9;
		16'h6766: out_word = 8'h4F;
		16'h6767: out_word = 8'h2E;
		16'h6768: out_word = 8'h4B;
		16'h6769: out_word = 8'h2E;
		16'h676A: out_word = 8'h00;
		16'h676B: out_word = 8'h56;
		16'h676C: out_word = 8'h65;
		16'h676D: out_word = 8'h72;
		16'h676E: out_word = 8'h69;
		16'h676F: out_word = 8'h66;
		16'h6770: out_word = 8'h79;
		16'h6771: out_word = 8'h20;
		16'h6772: out_word = 8'h45;
		16'h6773: out_word = 8'h72;
		16'h6774: out_word = 8'h72;
		16'h6775: out_word = 8'h6F;
		16'h6776: out_word = 8'h72;
		16'h6777: out_word = 8'h2E;
		16'h6778: out_word = 8'h8D;
		16'h6779: out_word = 8'h42;
		16'h677A: out_word = 8'h41;
		16'h677B: out_word = 8'h43;
		16'h677C: out_word = 8'h4B;
		16'h677D: out_word = 8'h55;
		16'h677E: out_word = 8'h50;
		16'h677F: out_word = 8'h20;
		16'h6780: out_word = 8'h44;
		16'h6781: out_word = 8'h49;
		16'h6782: out_word = 8'h53;
		16'h6783: out_word = 8'h4B;
		16'h6784: out_word = 8'h8D;
		16'h6785: out_word = 8'h49;
		16'h6786: out_word = 8'h6E;
		16'h6787: out_word = 8'h73;
		16'h6788: out_word = 8'h65;
		16'h6789: out_word = 8'h72;
		16'h678A: out_word = 8'h74;
		16'h678B: out_word = 8'h20;
		16'h678C: out_word = 8'h44;
		16'h678D: out_word = 8'h65;
		16'h678E: out_word = 8'h73;
		16'h678F: out_word = 8'h74;
		16'h6790: out_word = 8'h69;
		16'h6791: out_word = 8'h6E;
		16'h6792: out_word = 8'h61;
		16'h6793: out_word = 8'h74;
		16'h6794: out_word = 8'h69;
		16'h6795: out_word = 8'h6F;
		16'h6796: out_word = 8'h6E;
		16'h6797: out_word = 8'h20;
		16'h6798: out_word = 8'h64;
		16'h6799: out_word = 8'h69;
		16'h679A: out_word = 8'h73;
		16'h679B: out_word = 8'h6B;
		16'h679C: out_word = 8'h0D;
		16'h679D: out_word = 8'h74;
		16'h679E: out_word = 8'h68;
		16'h679F: out_word = 8'h65;
		16'h67A0: out_word = 8'h6E;
		16'h67A1: out_word = 8'h20;
		16'h67A2: out_word = 8'h70;
		16'h67A3: out_word = 8'h72;
		16'h67A4: out_word = 8'h65;
		16'h67A5: out_word = 8'h73;
		16'h67A6: out_word = 8'h73;
		16'h67A7: out_word = 8'h20;
		16'h67A8: out_word = 8'h59;
		16'h67A9: out_word = 8'h00;
		16'h67AA: out_word = 8'h49;
		16'h67AB: out_word = 8'h6E;
		16'h67AC: out_word = 8'h73;
		16'h67AD: out_word = 8'h65;
		16'h67AE: out_word = 8'h72;
		16'h67AF: out_word = 8'h74;
		16'h67B0: out_word = 8'h20;
		16'h67B1: out_word = 8'h53;
		16'h67B2: out_word = 8'h6F;
		16'h67B3: out_word = 8'h75;
		16'h67B4: out_word = 8'h72;
		16'h67B5: out_word = 8'h63;
		16'h67B6: out_word = 8'h65;
		16'h67B7: out_word = 8'h20;
		16'h67B8: out_word = 8'h64;
		16'h67B9: out_word = 8'h69;
		16'h67BA: out_word = 8'h73;
		16'h67BB: out_word = 8'h6B;
		16'h67BC: out_word = 8'h20;
		16'h67BD: out_word = 8'h74;
		16'h67BE: out_word = 8'h68;
		16'h67BF: out_word = 8'h65;
		16'h67C0: out_word = 8'h6E;
		16'h67C1: out_word = 8'h20;
		16'h67C2: out_word = 8'h70;
		16'h67C3: out_word = 8'h72;
		16'h67C4: out_word = 8'h65;
		16'h67C5: out_word = 8'h73;
		16'h67C6: out_word = 8'h73;
		16'h67C7: out_word = 8'h20;
		16'h67C8: out_word = 8'h59;
		16'h67C9: out_word = 8'h00;
		16'h67CA: out_word = 8'h2A;
		16'h67CB: out_word = 8'h42;
		16'h67CC: out_word = 8'h52;
		16'h67CD: out_word = 8'h45;
		16'h67CE: out_word = 8'h41;
		16'h67CF: out_word = 8'h4B;
		16'h67D0: out_word = 8'h2A;
		16'h67D1: out_word = 8'h8D;
		16'h67D2: out_word = 8'h4F;
		16'h67D3: out_word = 8'h75;
		16'h67D4: out_word = 8'h74;
		16'h67D5: out_word = 8'h20;
		16'h67D6: out_word = 8'h6F;
		16'h67D7: out_word = 8'h66;
		16'h67D8: out_word = 8'h20;
		16'h67D9: out_word = 8'h52;
		16'h67DA: out_word = 8'h41;
		16'h67DB: out_word = 8'h4D;
		16'h67DC: out_word = 8'h8D;
		16'h67DD: out_word = 8'h41;
		16'h67DE: out_word = 8'h72;
		16'h67DF: out_word = 8'h72;
		16'h67E0: out_word = 8'h61;
		16'h67E1: out_word = 8'h79;
		16'h67E2: out_word = 8'h20;
		16'h67E3: out_word = 8'h6E;
		16'h67E4: out_word = 8'h6F;
		16'h67E5: out_word = 8'h74;
		16'h67E6: out_word = 8'h20;
		16'h67E7: out_word = 8'h66;
		16'h67E8: out_word = 8'h6F;
		16'h67E9: out_word = 8'h75;
		16'h67EA: out_word = 8'h6E;
		16'h67EB: out_word = 8'h64;
		16'h67EC: out_word = 8'h8D;
		16'h67ED: out_word = 8'h44;
		16'h67EE: out_word = 8'h69;
		16'h67EF: out_word = 8'h72;
		16'h67F0: out_word = 8'h65;
		16'h67F1: out_word = 8'h63;
		16'h67F2: out_word = 8'h74;
		16'h67F3: out_word = 8'h6F;
		16'h67F4: out_word = 8'h72;
		16'h67F5: out_word = 8'h79;
		16'h67F6: out_word = 8'h20;
		16'h67F7: out_word = 8'h66;
		16'h67F8: out_word = 8'h75;
		16'h67F9: out_word = 8'h6C;
		16'h67FA: out_word = 8'h6C;
		16'h67FB: out_word = 8'h8D;
		16'h67FC: out_word = 8'h4E;
		16'h67FD: out_word = 8'h6F;
		16'h67FE: out_word = 8'h20;
		16'h67FF: out_word = 8'h64;
		16'h6800: out_word = 8'h69;
		16'h6801: out_word = 8'h73;
		16'h6802: out_word = 8'h6B;
		16'h6803: out_word = 8'h8D;
		16'h6804: out_word = 8'h53;
		16'h6805: out_word = 8'h74;
		16'h6806: out_word = 8'h72;
		16'h6807: out_word = 8'h65;
		16'h6808: out_word = 8'h61;
		16'h6809: out_word = 8'h6D;
		16'h680A: out_word = 8'h20;
		16'h680B: out_word = 8'h6F;
		16'h680C: out_word = 8'h70;
		16'h680D: out_word = 8'h65;
		16'h680E: out_word = 8'h6E;
		16'h680F: out_word = 8'h65;
		16'h6810: out_word = 8'h64;
		16'h6811: out_word = 8'h8D;
		16'h6812: out_word = 8'h4E;
		16'h6813: out_word = 8'h6F;
		16'h6814: out_word = 8'h74;
		16'h6815: out_word = 8'h20;
		16'h6816: out_word = 8'h64;
		16'h6817: out_word = 8'h69;
		16'h6818: out_word = 8'h73;
		16'h6819: out_word = 8'h6B;
		16'h681A: out_word = 8'h20;
		16'h681B: out_word = 8'h66;
		16'h681C: out_word = 8'h69;
		16'h681D: out_word = 8'h6C;
		16'h681E: out_word = 8'h65;
		16'h681F: out_word = 8'h8D;
		16'h6820: out_word = 8'h46;
		16'h6821: out_word = 8'h69;
		16'h6822: out_word = 8'h6C;
		16'h6823: out_word = 8'h65;
		16'h6824: out_word = 8'h20;
		16'h6825: out_word = 8'h65;
		16'h6826: out_word = 8'h78;
		16'h6827: out_word = 8'h69;
		16'h6828: out_word = 8'h73;
		16'h6829: out_word = 8'h74;
		16'h682A: out_word = 8'h73;
		16'h682B: out_word = 8'h0D;
		16'h682C: out_word = 8'h4F;
		16'h682D: out_word = 8'h76;
		16'h682E: out_word = 8'h65;
		16'h682F: out_word = 8'h72;
		16'h6830: out_word = 8'h20;
		16'h6831: out_word = 8'h77;
		16'h6832: out_word = 8'h72;
		16'h6833: out_word = 8'h69;
		16'h6834: out_word = 8'h74;
		16'h6835: out_word = 8'h65;
		16'h6836: out_word = 8'h3F;
		16'h6837: out_word = 8'h28;
		16'h6838: out_word = 8'h59;
		16'h6839: out_word = 8'h2F;
		16'h683A: out_word = 8'h4E;
		16'h683B: out_word = 8'hA9;
		16'h683C: out_word = 8'hF5;
		16'h683D: out_word = 8'hC5;
		16'h683E: out_word = 8'hED;
		16'h683F: out_word = 8'h53;
		16'h6840: out_word = 8'h04;
		16'h6841: out_word = 8'h5D;
		16'h6842: out_word = 8'h22;
		16'h6843: out_word = 8'h02;
		16'h6844: out_word = 8'h5D;
		16'h6845: out_word = 8'hCD;
		16'h6846: out_word = 8'hF1;
		16'h6847: out_word = 8'h20;
		16'h6848: out_word = 8'h3E;
		16'h6849: out_word = 8'hFF;
		16'h684A: out_word = 8'h32;
		16'h684B: out_word = 8'h15;
		16'h684C: out_word = 8'h5D;
		16'h684D: out_word = 8'h32;
		16'h684E: out_word = 8'h1F;
		16'h684F: out_word = 8'h5D;
		16'h6850: out_word = 8'hC1;
		16'h6851: out_word = 8'hF1;
		16'h6852: out_word = 8'h21;
		16'h6853: out_word = 8'h01;
		16'h6854: out_word = 8'h02;
		16'h6855: out_word = 8'h22;
		16'h6856: out_word = 8'h1A;
		16'h6857: out_word = 8'h5D;
		16'h6858: out_word = 8'h21;
		16'h6859: out_word = 8'h00;
		16'h685A: out_word = 8'h00;
		16'h685B: out_word = 8'h39;
		16'h685C: out_word = 8'h22;
		16'h685D: out_word = 8'h1C;
		16'h685E: out_word = 8'h5D;
		16'h685F: out_word = 8'h2B;
		16'h6860: out_word = 8'h2B;
		16'h6861: out_word = 8'hF9;
		16'h6862: out_word = 8'hF5;
		16'h6863: out_word = 8'hCD;
		16'h6864: out_word = 8'h1D;
		16'h6865: out_word = 8'h02;
		16'h6866: out_word = 8'h21;
		16'h6867: out_word = 8'h8C;
		16'h6868: out_word = 8'h28;
		16'h6869: out_word = 8'h7E;
		16'h686A: out_word = 8'hB9;
		16'h686B: out_word = 8'h20;
		16'h686C: out_word = 8'h12;
		16'h686D: out_word = 8'hF1;
		16'h686E: out_word = 8'h23;
		16'h686F: out_word = 8'h5E;
		16'h6870: out_word = 8'h23;
		16'h6871: out_word = 8'h56;
		16'h6872: out_word = 8'h21;
		16'h6873: out_word = 8'hD3;
		16'h6874: out_word = 8'h01;
		16'h6875: out_word = 8'hE5;
		16'h6876: out_word = 8'hD5;
		16'h6877: out_word = 8'h2A;
		16'h6878: out_word = 8'h02;
		16'h6879: out_word = 8'h5D;
		16'h687A: out_word = 8'hED;
		16'h687B: out_word = 8'h5B;
		16'h687C: out_word = 8'h04;
		16'h687D: out_word = 8'h5D;
		16'h687E: out_word = 8'hC9;
		16'h687F: out_word = 8'hFE;
		16'h6880: out_word = 8'hFF;
		16'h6881: out_word = 8'h20;
		16'h6882: out_word = 8'h04;
		16'h6883: out_word = 8'hF1;
		16'h6884: out_word = 8'hC3;
		16'h6885: out_word = 8'hD3;
		16'h6886: out_word = 8'h01;
		16'h6887: out_word = 8'h23;
		16'h6888: out_word = 8'h23;
		16'h6889: out_word = 8'h23;
		16'h688A: out_word = 8'h18;
		16'h688B: out_word = 8'hDD;
		16'h688C: out_word = 8'h00;
		16'h688D: out_word = 8'h98;
		16'h688E: out_word = 8'h3D;
		16'h688F: out_word = 8'h01;
		16'h6890: out_word = 8'hCB;
		16'h6891: out_word = 8'h3D;
		16'h6892: out_word = 8'h02;
		16'h6893: out_word = 8'h63;
		16'h6894: out_word = 8'h3E;
		16'h6895: out_word = 8'h03;
		16'h6896: out_word = 8'h02;
		16'h6897: out_word = 8'h3F;
		16'h6898: out_word = 8'h04;
		16'h6899: out_word = 8'h06;
		16'h689A: out_word = 8'h3F;
		16'h689B: out_word = 8'h05;
		16'h689C: out_word = 8'h3D;
		16'h689D: out_word = 8'h1E;
		16'h689E: out_word = 8'h06;
		16'h689F: out_word = 8'h4D;
		16'h68A0: out_word = 8'h1E;
		16'h68A1: out_word = 8'h07;
		16'h68A2: out_word = 8'hD8;
		16'h68A3: out_word = 8'h28;
		16'h68A4: out_word = 8'h08;
		16'h68A5: out_word = 8'h5C;
		16'h68A6: out_word = 8'h16;
		16'h68A7: out_word = 8'h09;
		16'h68A8: out_word = 8'h64;
		16'h68A9: out_word = 8'h16;
		16'h68AA: out_word = 8'h0A;
		16'h68AB: out_word = 8'hF0;
		16'h68AC: out_word = 8'h1C;
		16'h68AD: out_word = 8'h0B;
		16'h68AE: out_word = 8'hFB;
		16'h68AF: out_word = 8'h28;
		16'h68B0: out_word = 8'h0C;
		16'h68B1: out_word = 8'hF2;
		16'h68B2: out_word = 8'h28;
		16'h68B3: out_word = 8'h0D;
		16'h68B4: out_word = 8'h10;
		16'h68B5: out_word = 8'h3C;
		16'h68B6: out_word = 8'h0E;
		16'h68B7: out_word = 8'h0F;
		16'h68B8: out_word = 8'h29;
		16'h68B9: out_word = 8'h0F;
		16'h68BA: out_word = 8'h14;
		16'h68BB: out_word = 8'h3C;
		16'h68BC: out_word = 8'h10;
		16'h68BD: out_word = 8'h18;
		16'h68BE: out_word = 8'h3C;
		16'h68BF: out_word = 8'h11;
		16'h68C0: out_word = 8'h1D;
		16'h68C1: out_word = 8'h3C;
		16'h68C2: out_word = 8'h12;
		16'h68C3: out_word = 8'h26;
		16'h68C4: out_word = 8'h29;
		16'h68C5: out_word = 8'h13;
		16'h68C6: out_word = 8'hE0;
		16'h68C7: out_word = 8'h28;
		16'h68C8: out_word = 8'h14;
		16'h68C9: out_word = 8'hE3;
		16'h68CA: out_word = 8'h28;
		16'h68CB: out_word = 8'h15;
		16'h68CC: out_word = 8'h39;
		16'h68CD: out_word = 8'h27;
		16'h68CE: out_word = 8'h16;
		16'h68CF: out_word = 8'hEB;
		16'h68D0: out_word = 8'h1F;
		16'h68D1: out_word = 8'h17;
		16'h68D2: out_word = 8'hF6;
		16'h68D3: out_word = 8'h1F;
		16'h68D4: out_word = 8'h18;
		16'h68D5: out_word = 8'h05;
		16'h68D6: out_word = 8'h04;
		16'h68D7: out_word = 8'hFF;
		16'h68D8: out_word = 8'hF5;
		16'h68D9: out_word = 8'hCD;
		16'h68DA: out_word = 8'h05;
		16'h68DB: out_word = 8'h04;
		16'h68DC: out_word = 8'hF1;
		16'h68DD: out_word = 8'hC3;
		16'h68DE: out_word = 8'h79;
		16'h68DF: out_word = 8'h04;
		16'h68E0: out_word = 8'hAF;
		16'h68E1: out_word = 8'h18;
		16'h68E2: out_word = 8'h02;
		16'h68E3: out_word = 8'h3E;
		16'h68E4: out_word = 8'hFF;
		16'h68E5: out_word = 8'h11;
		16'h68E6: out_word = 8'hDD;
		16'h68E7: out_word = 8'h5C;
		16'h68E8: out_word = 8'h01;
		16'h68E9: out_word = 8'h10;
		16'h68EA: out_word = 8'h00;
		16'h68EB: out_word = 8'hB7;
		16'h68EC: out_word = 8'h28;
		16'h68ED: out_word = 8'h01;
		16'h68EE: out_word = 8'hEB;
		16'h68EF: out_word = 8'hED;
		16'h68F0: out_word = 8'hB0;
		16'h68F1: out_word = 8'hC9;
		16'h68F2: out_word = 8'hCD;
		16'h68F3: out_word = 8'h05;
		16'h68F4: out_word = 8'h04;
		16'h68F5: out_word = 8'hCD;
		16'h68F6: out_word = 8'hC4;
		16'h68F7: out_word = 8'h1A;
		16'h68F8: out_word = 8'hC3;
		16'h68F9: out_word = 8'h27;
		16'h68FA: out_word = 8'h1B;
		16'h68FB: out_word = 8'h22;
		16'h68FC: out_word = 8'hD7;
		16'h68FD: out_word = 8'h5C;
		16'h68FE: out_word = 8'hED;
		16'h68FF: out_word = 8'h53;
		16'h6900: out_word = 8'hD9;
		16'h6901: out_word = 8'h5C;
		16'h6902: out_word = 8'hED;
		16'h6903: out_word = 8'h53;
		16'h6904: out_word = 8'hDB;
		16'h6905: out_word = 8'h5C;
		16'h6906: out_word = 8'hC3;
		16'h6907: out_word = 8'hE6;
		16'h6908: out_word = 8'h33;
		16'h6909: out_word = 8'hCD;
		16'h690A: out_word = 8'hC4;
		16'h690B: out_word = 8'h1A;
		16'h690C: out_word = 8'hC3;
		16'h690D: out_word = 8'h71;
		16'h690E: out_word = 8'h33;
		16'h690F: out_word = 8'hB7;
		16'h6910: out_word = 8'h32;
		16'h6911: out_word = 8'hD6;
		16'h6912: out_word = 8'h5C;
		16'h6913: out_word = 8'h22;
		16'h6914: out_word = 8'hD9;
		16'h6915: out_word = 8'h5C;
		16'h6916: out_word = 8'hED;
		16'h6917: out_word = 8'h53;
		16'h6918: out_word = 8'hDB;
		16'h6919: out_word = 8'h5C;
		16'h691A: out_word = 8'hCD;
		16'h691B: out_word = 8'hB3;
		16'h691C: out_word = 8'h1C;
		16'h691D: out_word = 8'hCD;
		16'h691E: out_word = 8'hA4;
		16'h691F: out_word = 8'h18;
		16'h6920: out_word = 8'hCD;
		16'h6921: out_word = 8'hAB;
		16'h6922: out_word = 8'h18;
		16'h6923: out_word = 8'hC3;
		16'h6924: out_word = 8'h21;
		16'h6925: out_word = 8'h19;
		16'h6926: out_word = 8'hCD;
		16'h6927: out_word = 8'h05;
		16'h6928: out_word = 8'h04;
		16'h6929: out_word = 8'hCD;
		16'h692A: out_word = 8'hB3;
		16'h692B: out_word = 8'h1C;
		16'h692C: out_word = 8'hC3;
		16'h692D: out_word = 8'hA0;
		16'h692E: out_word = 8'h07;
		16'h692F: out_word = 8'hCD;
		16'h6930: out_word = 8'h57;
		16'h6931: out_word = 8'h1C;
		16'h6932: out_word = 8'hCD;
		16'h6933: out_word = 8'h05;
		16'h6934: out_word = 8'h04;
		16'h6935: out_word = 8'hC3;
		16'h6936: out_word = 8'hB3;
		16'h6937: out_word = 8'h1C;
		16'h6938: out_word = 8'hC5;
		16'h6939: out_word = 8'h06;
		16'h693A: out_word = 8'h08;
		16'h693B: out_word = 8'h7E;
		16'h693C: out_word = 8'hD7;
		16'h693D: out_word = 8'h23;
		16'h693E: out_word = 8'h10;
		16'h693F: out_word = 8'hFB;
		16'h6940: out_word = 8'h3E;
		16'h6941: out_word = 8'h3C;
		16'h6942: out_word = 8'hD7;
		16'h6943: out_word = 8'h7E;
		16'h6944: out_word = 8'hD7;
		16'h6945: out_word = 8'h3E;
		16'h6946: out_word = 8'h3E;
		16'h6947: out_word = 8'hD7;
		16'h6948: out_word = 8'hC1;
		16'h6949: out_word = 8'hC9;
		16'h694A: out_word = 8'hE5;
		16'h694B: out_word = 8'hD5;
		16'h694C: out_word = 8'hC5;
		16'h694D: out_word = 8'hF5;
		16'h694E: out_word = 8'h21;
		16'h694F: out_word = 8'h0C;
		16'h6950: out_word = 8'h5D;
		16'h6951: out_word = 8'h7E;
		16'h6952: out_word = 8'hB7;
		16'h6953: out_word = 8'h28;
		16'h6954: out_word = 8'h3D;
		16'h6955: out_word = 8'hE5;
		16'h6956: out_word = 8'h01;
		16'h6957: out_word = 8'h01;
		16'h6958: out_word = 8'h01;
		16'h6959: out_word = 8'hC5;
		16'h695A: out_word = 8'hCD;
		16'h695B: out_word = 8'hFD;
		16'h695C: out_word = 8'h19;
		16'h695D: out_word = 8'hC1;
		16'h695E: out_word = 8'hE1;
		16'h695F: out_word = 8'h36;
		16'h6960: out_word = 8'h00;
		16'h6961: out_word = 8'h21;
		16'h6962: out_word = 8'h25;
		16'h6963: out_word = 8'h5D;
		16'h6964: out_word = 8'hCD;
		16'h6965: out_word = 8'h32;
		16'h6966: out_word = 8'h1E;
		16'h6967: out_word = 8'h2A;
		16'h6968: out_word = 8'h11;
		16'h6969: out_word = 8'h5D;
		16'h696A: out_word = 8'h01;
		16'h696B: out_word = 8'h01;
		16'h696C: out_word = 8'h01;
		16'h696D: out_word = 8'h09;
		16'h696E: out_word = 8'h18;
		16'h696F: out_word = 8'h1F;
		16'h6970: out_word = 8'hE5;
		16'h6971: out_word = 8'hD5;
		16'h6972: out_word = 8'hC5;
		16'h6973: out_word = 8'hF5;
		16'h6974: out_word = 8'h21;
		16'h6975: out_word = 8'h0C;
		16'h6976: out_word = 8'h5D;
		16'h6977: out_word = 8'h7E;
		16'h6978: out_word = 8'hB7;
		16'h6979: out_word = 8'h20;
		16'h697A: out_word = 8'h17;
		16'h697B: out_word = 8'h36;
		16'h697C: out_word = 8'hFF;
		16'h697D: out_word = 8'h21;
		16'h697E: out_word = 8'h25;
		16'h697F: out_word = 8'h5D;
		16'h6980: out_word = 8'h01;
		16'h6981: out_word = 8'h01;
		16'h6982: out_word = 8'h01;
		16'h6983: out_word = 8'hCD;
		16'h6984: out_word = 8'h2E;
		16'h6985: out_word = 8'h1E;
		16'h6986: out_word = 8'hB7;
		16'h6987: out_word = 8'h01;
		16'h6988: out_word = 8'h01;
		16'h6989: out_word = 8'h01;
		16'h698A: out_word = 8'h2A;
		16'h698B: out_word = 8'h11;
		16'h698C: out_word = 8'h5D;
		16'h698D: out_word = 8'hED;
		16'h698E: out_word = 8'h42;
		16'h698F: out_word = 8'h22;
		16'h6990: out_word = 8'h11;
		16'h6991: out_word = 8'h5D;
		16'h6992: out_word = 8'hF1;
		16'h6993: out_word = 8'hC1;
		16'h6994: out_word = 8'hD1;
		16'h6995: out_word = 8'hE1;
		16'h6996: out_word = 8'hC9;
		16'h6997: out_word = 8'hAF;
		16'h6998: out_word = 8'h32;
		16'h6999: out_word = 8'hD7;
		16'h699A: out_word = 8'h5C;
		16'h699B: out_word = 8'hCD;
		16'h699C: out_word = 8'h75;
		16'h699D: out_word = 8'h1D;
		16'h699E: out_word = 8'hCD;
		16'h699F: out_word = 8'h2B;
		16'h69A0: out_word = 8'h04;
		16'h69A1: out_word = 8'hCA;
		16'h69A2: out_word = 8'h1A;
		16'h69A3: out_word = 8'h1D;
		16'h69A4: out_word = 8'hCD;
		16'h69A5: out_word = 8'h11;
		16'h69A6: out_word = 8'h3E;
		16'h69A7: out_word = 8'h3A;
		16'h69A8: out_word = 8'hD7;
		16'h69A9: out_word = 8'h5C;
		16'h69AA: out_word = 8'h77;
		16'h69AB: out_word = 8'hC3;
		16'h69AC: out_word = 8'hE1;
		16'h69AD: out_word = 8'h03;
		16'h69AE: out_word = 8'h3E;
		16'h69AF: out_word = 8'h80;
		16'h69B0: out_word = 8'h18;
		16'h69B1: out_word = 8'hE6;
		16'h69B2: out_word = 8'h0D;
		16'h69B3: out_word = 8'h2A;
		16'h69B4: out_word = 8'h45;
		16'h69B5: out_word = 8'h52;
		16'h69B6: out_word = 8'h52;
		16'h69B7: out_word = 8'h4F;
		16'h69B8: out_word = 8'h52;
		16'h69B9: out_word = 8'h2A;
		16'h69BA: out_word = 8'h8D;
		16'h69BB: out_word = 8'h0D;
		16'h69BC: out_word = 8'h4E;
		16'h69BD: out_word = 8'h6F;
		16'h69BE: out_word = 8'h20;
		16'h69BF: out_word = 8'h73;
		16'h69C0: out_word = 8'h70;
		16'h69C1: out_word = 8'h61;
		16'h69C2: out_word = 8'h63;
		16'h69C3: out_word = 8'h65;
		16'h69C4: out_word = 8'h8D;
		16'h69C5: out_word = 8'h0D;
		16'h69C6: out_word = 8'h46;
		16'h69C7: out_word = 8'h69;
		16'h69C8: out_word = 8'h6C;
		16'h69C9: out_word = 8'h65;
		16'h69CA: out_word = 8'h20;
		16'h69CB: out_word = 8'h65;
		16'h69CC: out_word = 8'h78;
		16'h69CD: out_word = 8'h69;
		16'h69CE: out_word = 8'h73;
		16'h69CF: out_word = 8'h74;
		16'h69D0: out_word = 8'h73;
		16'h69D1: out_word = 8'h8D;
		16'h69D2: out_word = 8'h20;
		16'h69D3: out_word = 8'h46;
		16'h69D4: out_word = 8'h72;
		16'h69D5: out_word = 8'h65;
		16'h69D6: out_word = 8'h65;
		16'h69D7: out_word = 8'h8D;
		16'h69D8: out_word = 8'h0D;
		16'h69D9: out_word = 8'h52;
		16'h69DA: out_word = 8'h65;
		16'h69DB: out_word = 8'h61;
		16'h69DC: out_word = 8'h64;
		16'h69DD: out_word = 8'h20;
		16'h69DE: out_word = 8'h4F;
		16'h69DF: out_word = 8'h6E;
		16'h69E0: out_word = 8'h6C;
		16'h69E1: out_word = 8'hF9;
		16'h69E2: out_word = 8'h0D;
		16'h69E3: out_word = 8'h44;
		16'h69E4: out_word = 8'h69;
		16'h69E5: out_word = 8'h73;
		16'h69E6: out_word = 8'h6B;
		16'h69E7: out_word = 8'h20;
		16'h69E8: out_word = 8'h45;
		16'h69E9: out_word = 8'h72;
		16'h69EA: out_word = 8'h72;
		16'h69EB: out_word = 8'h6F;
		16'h69EC: out_word = 8'hF2;
		16'h69ED: out_word = 8'h0D;
		16'h69EE: out_word = 8'h52;
		16'h69EF: out_word = 8'h65;
		16'h69F0: out_word = 8'h63;
		16'h69F1: out_word = 8'h2E;
		16'h69F2: out_word = 8'h20;
		16'h69F3: out_word = 8'h20;
		16'h69F4: out_word = 8'h4F;
		16'h69F5: out_word = 8'h2F;
		16'h69F6: out_word = 8'hC6;
		16'h69F7: out_word = 8'h54;
		16'h69F8: out_word = 8'h69;
		16'h69F9: out_word = 8'h74;
		16'h69FA: out_word = 8'h6C;
		16'h69FB: out_word = 8'h65;
		16'h69FC: out_word = 8'h3A;
		16'h69FD: out_word = 8'hA0;
		16'h69FE: out_word = 8'h0D;
		16'h69FF: out_word = 8'h52;
		16'h6A00: out_word = 8'h65;
		16'h6A01: out_word = 8'h74;
		16'h6A02: out_word = 8'h72;
		16'h6A03: out_word = 8'h79;
		16'h6A04: out_word = 8'h2C;
		16'h6A05: out_word = 8'h41;
		16'h6A06: out_word = 8'h62;
		16'h6A07: out_word = 8'h6F;
		16'h6A08: out_word = 8'h72;
		16'h6A09: out_word = 8'h74;
		16'h6A0A: out_word = 8'h2C;
		16'h6A0B: out_word = 8'h49;
		16'h6A0C: out_word = 8'h67;
		16'h6A0D: out_word = 8'h6E;
		16'h6A0E: out_word = 8'h6F;
		16'h6A0F: out_word = 8'h72;
		16'h6A10: out_word = 8'h65;
		16'h6A11: out_word = 8'h3F;
		16'h6A12: out_word = 8'h00;
		16'h6A13: out_word = 8'h0D;
		16'h6A14: out_word = 8'h54;
		16'h6A15: out_word = 8'h72;
		16'h6A16: out_word = 8'h6B;
		16'h6A17: out_word = 8'hA0;
		16'h6A18: out_word = 8'h20;
		16'h6A19: out_word = 8'h73;
		16'h6A1A: out_word = 8'h65;
		16'h6A1B: out_word = 8'h63;
		16'h6A1C: out_word = 8'hA0;
		16'h6A1D: out_word = 8'h20;
		16'h6A1E: out_word = 8'h44;
		16'h6A1F: out_word = 8'h65;
		16'h6A20: out_word = 8'h6C;
		16'h6A21: out_word = 8'h2E;
		16'h6A22: out_word = 8'h20;
		16'h6A23: out_word = 8'h46;
		16'h6A24: out_word = 8'h69;
		16'h6A25: out_word = 8'h6C;
		16'h6A26: out_word = 8'h65;
		16'h6A27: out_word = 8'h8D;
		16'h6A28: out_word = 8'h0D;
		16'h6A29: out_word = 8'h4E;
		16'h6A2A: out_word = 8'h6F;
		16'h6A2B: out_word = 8'h20;
		16'h6A2C: out_word = 8'h46;
		16'h6A2D: out_word = 8'h69;
		16'h6A2E: out_word = 8'h6C;
		16'h6A2F: out_word = 8'h65;
		16'h6A30: out_word = 8'h28;
		16'h6A31: out_word = 8'h73;
		16'h6A32: out_word = 8'h29;
		16'h6A33: out_word = 8'h8D;
		16'h6A34: out_word = 8'h00;
		16'h6A35: out_word = 8'h21;
		16'h6A36: out_word = 8'h41;
		16'h6A37: out_word = 8'h2A;
		16'h6A38: out_word = 8'h11;
		16'h6A39: out_word = 8'h80;
		16'h6A3A: out_word = 8'h40;
		16'h6A3B: out_word = 8'h01;
		16'h6A3C: out_word = 8'h20;
		16'h6A3D: out_word = 8'h00;
		16'h6A3E: out_word = 8'hED;
		16'h6A3F: out_word = 8'hB0;
		16'h6A40: out_word = 8'hC9;
		16'h6A41: out_word = 8'h3A;
		16'h6A42: out_word = 8'hB5;
		16'h6A43: out_word = 8'h03;
		16'h6A44: out_word = 8'hFE;
		16'h6A45: out_word = 8'hF3;
		16'h6A46: out_word = 8'h3E;
		16'h6A47: out_word = 8'h10;
		16'h6A48: out_word = 8'h28;
		16'h6A49: out_word = 8'h01;
		16'h6A4A: out_word = 8'hAF;
		16'h6A4B: out_word = 8'h32;
		16'h6A4C: out_word = 8'h01;
		16'h6A4D: out_word = 8'h5C;
		16'h6A4E: out_word = 8'h01;
		16'h6A4F: out_word = 8'hFD;
		16'h6A50: out_word = 8'h7F;
		16'h6A51: out_word = 8'h3E;
		16'h6A52: out_word = 8'h10;
		16'h6A53: out_word = 8'hED;
		16'h6A54: out_word = 8'h79;
		16'h6A55: out_word = 8'hC9;
		16'h6A56: out_word = 8'hC3;
		16'h6A57: out_word = 8'h1A;
		16'h6A58: out_word = 8'h0A;
		16'h6A59: out_word = 8'hE5;
		16'h6A5A: out_word = 8'hDD;
		16'h6A5B: out_word = 8'hE5;
		16'h6A5C: out_word = 8'hFD;
		16'h6A5D: out_word = 8'hE5;
		16'h6A5E: out_word = 8'hD9;
		16'h6A5F: out_word = 8'hC5;
		16'h6A60: out_word = 8'hD5;
		16'h6A61: out_word = 8'hE5;
		16'h6A62: out_word = 8'h08;
		16'h6A63: out_word = 8'hF5;
		16'h6A64: out_word = 8'hED;
		16'h6A65: out_word = 8'h57;
		16'h6A66: out_word = 8'hF5;
		16'h6A67: out_word = 8'hED;
		16'h6A68: out_word = 8'h5F;
		16'h6A69: out_word = 8'hF5;
		16'h6A6A: out_word = 8'h21;
		16'h6A6B: out_word = 8'h00;
		16'h6A6C: out_word = 8'h00;
		16'h6A6D: out_word = 8'h39;
		16'h6A6E: out_word = 8'hE5;
		16'h6A6F: out_word = 8'hCD;
		16'h6A70: out_word = 8'h01;
		16'h6A71: out_word = 8'h0A;
		16'h6A72: out_word = 8'h00;
		16'h6A73: out_word = 8'h3E;
		16'h6A74: out_word = 8'h3F;
		16'h6A75: out_word = 8'hED;
		16'h6A76: out_word = 8'h47;
		16'h6A77: out_word = 8'hDB;
		16'h6A78: out_word = 8'h1F;
		16'h6A79: out_word = 8'hE6;
		16'h6A7A: out_word = 8'h80;
		16'h6A7B: out_word = 8'h0F;
		16'h6A7C: out_word = 8'h0F;
		16'h6A7D: out_word = 8'h0F;
		16'h6A7E: out_word = 8'h32;
		16'h6A7F: out_word = 8'h01;
		16'h6A80: out_word = 8'h5C;
		16'h6A81: out_word = 8'hCD;
		16'h6A82: out_word = 8'h65;
		16'h6A83: out_word = 8'h2F;
		16'h6A84: out_word = 8'hCD;
		16'h6A85: out_word = 8'hA0;
		16'h6A86: out_word = 8'h3E;
		16'h6A87: out_word = 8'hCD;
		16'h6A88: out_word = 8'hA0;
		16'h6A89: out_word = 8'h3E;
		16'h6A8A: out_word = 8'h11;
		16'h6A8B: out_word = 8'h0A;
		16'h6A8C: out_word = 8'h00;
		16'h6A8D: out_word = 8'h21;
		16'h6A8E: out_word = 8'h00;
		16'h6A8F: out_word = 8'h40;
		16'h6A90: out_word = 8'hE5;
		16'h6A91: out_word = 8'hCD;
		16'h6A92: out_word = 8'h73;
		16'h6A93: out_word = 8'h2D;
		16'h6A94: out_word = 8'h21;
		16'h6A95: out_word = 8'h00;
		16'h6A96: out_word = 8'h41;
		16'h6A97: out_word = 8'h11;
		16'h6A98: out_word = 8'h0B;
		16'h6A99: out_word = 8'h00;
		16'h6A9A: out_word = 8'hCD;
		16'h6A9B: out_word = 8'h73;
		16'h6A9C: out_word = 8'h2D;
		16'h6A9D: out_word = 8'hE1;
		16'h6A9E: out_word = 8'hE5;
		16'h6A9F: out_word = 8'h11;
		16'h6AA0: out_word = 8'h08;
		16'h6AA1: out_word = 8'h00;
		16'h6AA2: out_word = 8'hCD;
		16'h6AA3: out_word = 8'h1B;
		16'h6AA4: out_word = 8'h2F;
		16'h6AA5: out_word = 8'h21;
		16'h6AA6: out_word = 8'hE3;
		16'h6AA7: out_word = 8'h40;
		16'h6AA8: out_word = 8'h7E;
		16'h6AA9: out_word = 8'h32;
		16'h6AAA: out_word = 8'h00;
		16'h6AAB: out_word = 8'h5C;
		16'h6AAC: out_word = 8'h23;
		16'h6AAD: out_word = 8'h7E;
		16'h6AAE: out_word = 8'h34;
		16'h6AAF: out_word = 8'h23;
		16'h6AB0: out_word = 8'h5E;
		16'h6AB1: out_word = 8'h23;
		16'h6AB2: out_word = 8'h56;
		16'h6AB3: out_word = 8'hB7;
		16'h6AB4: out_word = 8'hEB;
		16'h6AB5: out_word = 8'h11;
		16'h6AB6: out_word = 8'hC0;
		16'h6AB7: out_word = 8'h00;
		16'h6AB8: out_word = 8'hED;
		16'h6AB9: out_word = 8'h52;
		16'h6ABA: out_word = 8'h22;
		16'h6ABB: out_word = 8'hE5;
		16'h6ABC: out_word = 8'h40;
		16'h6ABD: out_word = 8'h21;
		16'h6ABE: out_word = 8'h00;
		16'h6ABF: out_word = 8'h40;
		16'h6AC0: out_word = 8'h11;
		16'h6AC1: out_word = 8'h08;
		16'h6AC2: out_word = 8'h00;
		16'h6AC3: out_word = 8'hCD;
		16'h6AC4: out_word = 8'h73;
		16'h6AC5: out_word = 8'h2D;
		16'h6AC6: out_word = 8'hE1;
		16'h6AC7: out_word = 8'hED;
		16'h6AC8: out_word = 8'h5B;
		16'h6AC9: out_word = 8'hE1;
		16'h6ACA: out_word = 8'h40;
		16'h6ACB: out_word = 8'hD5;
		16'h6ACC: out_word = 8'h11;
		16'h6ACD: out_word = 8'h0A;
		16'h6ACE: out_word = 8'h00;
		16'h6ACF: out_word = 8'hCD;
		16'h6AD0: out_word = 8'h1B;
		16'h6AD1: out_word = 8'h2F;
		16'h6AD2: out_word = 8'hD1;
		16'h6AD3: out_word = 8'hCD;
		16'h6AD4: out_word = 8'h4C;
		16'h6AD5: out_word = 8'h2D;
		16'h6AD6: out_word = 8'hD5;
		16'h6AD7: out_word = 8'h3E;
		16'h6AD8: out_word = 8'h3C;
		16'h6AD9: out_word = 8'hD3;
		16'h6ADA: out_word = 8'hFF;
		16'h6ADB: out_word = 8'hCD;
		16'h6ADC: out_word = 8'h65;
		16'h6ADD: out_word = 8'h2F;
		16'h6ADE: out_word = 8'h21;
		16'h6ADF: out_word = 8'h00;
		16'h6AE0: out_word = 8'h40;
		16'h6AE1: out_word = 8'h11;
		16'h6AE2: out_word = 8'h08;
		16'h6AE3: out_word = 8'h00;
		16'h6AE4: out_word = 8'h06;
		16'h6AE5: out_word = 8'h01;
		16'h6AE6: out_word = 8'hCD;
		16'h6AE7: out_word = 8'h1B;
		16'h6AE8: out_word = 8'h2F;
		16'h6AE9: out_word = 8'hD1;
		16'h6AEA: out_word = 8'h2A;
		16'h6AEB: out_word = 8'hE1;
		16'h6AEC: out_word = 8'h40;
		16'h6AED: out_word = 8'hED;
		16'h6AEE: out_word = 8'h53;
		16'h6AEF: out_word = 8'hE1;
		16'h6AF0: out_word = 8'h40;
		16'h6AF1: out_word = 8'hE5;
		16'h6AF2: out_word = 8'h21;
		16'h6AF3: out_word = 8'h00;
		16'h6AF4: out_word = 8'h40;
		16'h6AF5: out_word = 8'h11;
		16'h6AF6: out_word = 8'h08;
		16'h6AF7: out_word = 8'h00;
		16'h6AF8: out_word = 8'h06;
		16'h6AF9: out_word = 8'h01;
		16'h6AFA: out_word = 8'hCD;
		16'h6AFB: out_word = 8'h73;
		16'h6AFC: out_word = 8'h2D;
		16'h6AFD: out_word = 8'h3A;
		16'h6AFE: out_word = 8'hE4;
		16'h6AFF: out_word = 8'h40;
		16'h6B00: out_word = 8'h3D;
		16'h6B01: out_word = 8'hCD;
		16'h6B02: out_word = 8'hE5;
		16'h6B03: out_word = 8'h2C;
		16'h6B04: out_word = 8'h36;
		16'h6B05: out_word = 8'h40;
		16'h6B06: out_word = 8'h23;
		16'h6B07: out_word = 8'h06;
		16'h6B08: out_word = 8'h07;
		16'h6B09: out_word = 8'h36;
		16'h6B0A: out_word = 8'h20;
		16'h6B0B: out_word = 8'h23;
		16'h6B0C: out_word = 8'h10;
		16'h6B0D: out_word = 8'hFB;
		16'h6B0E: out_word = 8'h36;
		16'h6B0F: out_word = 8'h43;
		16'h6B10: out_word = 8'hD1;
		16'h6B11: out_word = 8'hC1;
		16'h6B12: out_word = 8'h23;
		16'h6B13: out_word = 8'h71;
		16'h6B14: out_word = 8'h23;
		16'h6B15: out_word = 8'h70;
		16'h6B16: out_word = 8'h23;
		16'h6B17: out_word = 8'h23;
		16'h6B18: out_word = 8'h23;
		16'h6B19: out_word = 8'h36;
		16'h6B1A: out_word = 8'hC0;
		16'h6B1B: out_word = 8'h23;
		16'h6B1C: out_word = 8'h73;
		16'h6B1D: out_word = 8'h23;
		16'h6B1E: out_word = 8'h72;
		16'h6B1F: out_word = 8'h21;
		16'h6B20: out_word = 8'h00;
		16'h6B21: out_word = 8'h40;
		16'h6B22: out_word = 8'h11;
		16'h6B23: out_word = 8'h00;
		16'h6B24: out_word = 8'h00;
		16'h6B25: out_word = 8'hDB;
		16'h6B26: out_word = 8'h5F;
		16'h6B27: out_word = 8'h3D;
		16'h6B28: out_word = 8'h5F;
		16'h6B29: out_word = 8'h06;
		16'h6B2A: out_word = 8'h01;
		16'h6B2B: out_word = 8'hCD;
		16'h6B2C: out_word = 8'h73;
		16'h6B2D: out_word = 8'h2D;
		16'h6B2E: out_word = 8'h21;
		16'h6B2F: out_word = 8'h00;
		16'h6B30: out_word = 8'h00;
		16'h6B31: out_word = 8'h39;
		16'h6B32: out_word = 8'h22;
		16'h6B33: out_word = 8'h40;
		16'h6B34: out_word = 8'h41;
		16'h6B35: out_word = 8'h31;
		16'h6B36: out_word = 8'hFF;
		16'h6B37: out_word = 8'h41;
		16'h6B38: out_word = 8'hCD;
		16'h6B39: out_word = 8'h35;
		16'h6B3A: out_word = 8'h2A;
		16'h6B3B: out_word = 8'h21;
		16'h6B3C: out_word = 8'h00;
		16'h6B3D: out_word = 8'hC0;
		16'h6B3E: out_word = 8'hAF;
		16'h6B3F: out_word = 8'h86;
		16'h6B40: out_word = 8'h23;
		16'h6B41: out_word = 8'h47;
		16'h6B42: out_word = 8'h7C;
		16'h6B43: out_word = 8'hB7;
		16'h6B44: out_word = 8'h78;
		16'h6B45: out_word = 8'h20;
		16'h6B46: out_word = 8'hF8;
		16'h6B47: out_word = 8'h21;
		16'h6B48: out_word = 8'h00;
		16'h6B49: out_word = 8'h41;
		16'h6B4A: out_word = 8'h77;
		16'h6B4B: out_word = 8'hE5;
		16'h6B4C: out_word = 8'h21;
		16'h6B4D: out_word = 8'h58;
		16'h6B4E: out_word = 8'h2B;
		16'h6B4F: out_word = 8'hE5;
		16'h6B50: out_word = 8'h21;
		16'h6B51: out_word = 8'h2F;
		16'h6B52: out_word = 8'h3D;
		16'h6B53: out_word = 8'hE5;
		16'h6B54: out_word = 8'hF3;
		16'h6B55: out_word = 8'hC3;
		16'h6B56: out_word = 8'h80;
		16'h6B57: out_word = 8'h40;
		16'h6B58: out_word = 8'hE1;
		16'h6B59: out_word = 8'h01;
		16'h6B5A: out_word = 8'hFD;
		16'h6B5B: out_word = 8'h7F;
		16'h6B5C: out_word = 8'h3E;
		16'h6B5D: out_word = 8'hAA;
		16'h6B5E: out_word = 8'h32;
		16'h6B5F: out_word = 8'h30;
		16'h6B60: out_word = 8'h41;
		16'h6B61: out_word = 8'h16;
		16'h6B62: out_word = 8'h05;
		16'h6B63: out_word = 8'h3A;
		16'h6B64: out_word = 8'h01;
		16'h6B65: out_word = 8'h5C;
		16'h6B66: out_word = 8'hB2;
		16'h6B67: out_word = 8'h57;
		16'h6B68: out_word = 8'hED;
		16'h6B69: out_word = 8'h51;
		16'h6B6A: out_word = 8'h3A;
		16'h6B6B: out_word = 8'h30;
		16'h6B6C: out_word = 8'hC1;
		16'h6B6D: out_word = 8'hFE;
		16'h6B6E: out_word = 8'hAA;
		16'h6B6F: out_word = 8'hC2;
		16'h6B70: out_word = 8'h1B;
		16'h6B71: out_word = 8'h2C;
		16'h6B72: out_word = 8'h7A;
		16'h6B73: out_word = 8'hE6;
		16'h6B74: out_word = 8'hF8;
		16'h6B75: out_word = 8'h57;
		16'h6B76: out_word = 8'h23;
		16'h6B77: out_word = 8'h72;
		16'h6B78: out_word = 8'hED;
		16'h6B79: out_word = 8'h51;
		16'h6B7A: out_word = 8'hAF;
		16'h6B7B: out_word = 8'h21;
		16'h6B7C: out_word = 8'h00;
		16'h6B7D: out_word = 8'hC0;
		16'h6B7E: out_word = 8'h86;
		16'h6B7F: out_word = 8'h23;
		16'h6B80: out_word = 8'h5F;
		16'h6B81: out_word = 8'h7C;
		16'h6B82: out_word = 8'hB7;
		16'h6B83: out_word = 8'h7B;
		16'h6B84: out_word = 8'h20;
		16'h6B85: out_word = 8'hF8;
		16'h6B86: out_word = 8'h21;
		16'h6B87: out_word = 8'h00;
		16'h6B88: out_word = 8'h41;
		16'h6B89: out_word = 8'hBE;
		16'h6B8A: out_word = 8'h23;
		16'h6B8B: out_word = 8'h28;
		16'h6B8C: out_word = 8'h06;
		16'h6B8D: out_word = 8'h14;
		16'h6B8E: out_word = 8'hCB;
		16'h6B8F: out_word = 8'h5A;
		16'h6B90: out_word = 8'h28;
		16'h6B91: out_word = 8'hE5;
		16'h6B92: out_word = 8'h15;
		16'h6B93: out_word = 8'h06;
		16'h6B94: out_word = 8'h08;
		16'h6B95: out_word = 8'hC5;
		16'h6B96: out_word = 8'hCD;
		16'h6B97: out_word = 8'h37;
		16'h6B98: out_word = 8'h2C;
		16'h6B99: out_word = 8'hC1;
		16'h6B9A: out_word = 8'h10;
		16'h6B9B: out_word = 8'hF9;
		16'h6B9C: out_word = 8'h0E;
		16'h6B9D: out_word = 8'h00;
		16'h6B9E: out_word = 8'hCD;
		16'h6B9F: out_word = 8'h3A;
		16'h6BA0: out_word = 8'h2F;
		16'h6BA1: out_word = 8'hCD;
		16'h6BA2: out_word = 8'h2A;
		16'h6BA3: out_word = 8'h2D;
		16'h6BA4: out_word = 8'h3A;
		16'h6BA5: out_word = 8'hE4;
		16'h6BA6: out_word = 8'h40;
		16'h6BA7: out_word = 8'h32;
		16'h6BA8: out_word = 8'h02;
		16'h6BA9: out_word = 8'h41;
		16'h6BAA: out_word = 8'h3C;
		16'h6BAB: out_word = 8'h32;
		16'h6BAC: out_word = 8'hE4;
		16'h6BAD: out_word = 8'h40;
		16'h6BAE: out_word = 8'h2A;
		16'h6BAF: out_word = 8'hE5;
		16'h6BB0: out_word = 8'h40;
		16'h6BB1: out_word = 8'h11;
		16'h6BB2: out_word = 8'h01;
		16'h6BB3: out_word = 8'h00;
		16'h6BB4: out_word = 8'hED;
		16'h6BB5: out_word = 8'h52;
		16'h6BB6: out_word = 8'h22;
		16'h6BB7: out_word = 8'hE5;
		16'h6BB8: out_word = 8'h40;
		16'h6BB9: out_word = 8'hD8;
		16'h6BBA: out_word = 8'h2A;
		16'h6BBB: out_word = 8'hE1;
		16'h6BBC: out_word = 8'h40;
		16'h6BBD: out_word = 8'h22;
		16'h6BBE: out_word = 8'h1E;
		16'h6BBF: out_word = 8'h41;
		16'h6BC0: out_word = 8'hCD;
		16'h6BC1: out_word = 8'h1E;
		16'h6BC2: out_word = 8'h2D;
		16'h6BC3: out_word = 8'h3E;
		16'h6BC4: out_word = 8'h38;
		16'h6BC5: out_word = 8'h32;
		16'h6BC6: out_word = 8'h11;
		16'h6BC7: out_word = 8'h41;
		16'h6BC8: out_word = 8'h3E;
		16'h6BC9: out_word = 8'h01;
		16'h6BCA: out_word = 8'h32;
		16'h6BCB: out_word = 8'h1D;
		16'h6BCC: out_word = 8'h41;
		16'h6BCD: out_word = 8'h21;
		16'h6BCE: out_word = 8'h00;
		16'h6BCF: out_word = 8'h41;
		16'h6BD0: out_word = 8'h22;
		16'h6BD1: out_word = 8'h19;
		16'h6BD2: out_word = 8'h41;
		16'h6BD3: out_word = 8'h21;
		16'h6BD4: out_word = 8'h00;
		16'h6BD5: out_word = 8'h01;
		16'h6BD6: out_word = 8'h22;
		16'h6BD7: out_word = 8'h1B;
		16'h6BD8: out_word = 8'h41;
		16'h6BD9: out_word = 8'hED;
		16'h6BDA: out_word = 8'h5B;
		16'h6BDB: out_word = 8'hE1;
		16'h6BDC: out_word = 8'h40;
		16'h6BDD: out_word = 8'hCD;
		16'h6BDE: out_word = 8'h65;
		16'h6BDF: out_word = 8'h2F;
		16'h6BE0: out_word = 8'h4A;
		16'h6BE1: out_word = 8'hCD;
		16'h6BE2: out_word = 8'h3A;
		16'h6BE3: out_word = 8'h2F;
		16'h6BE4: out_word = 8'h21;
		16'h6BE5: out_word = 8'h00;
		16'h6BE6: out_word = 8'h41;
		16'h6BE7: out_word = 8'h06;
		16'h6BE8: out_word = 8'h01;
		16'h6BE9: out_word = 8'hCD;
		16'h6BEA: out_word = 8'h58;
		16'h6BEB: out_word = 8'h2D;
		16'h6BEC: out_word = 8'hED;
		16'h6BED: out_word = 8'h53;
		16'h6BEE: out_word = 8'hE1;
		16'h6BEF: out_word = 8'h40;
		16'h6BF0: out_word = 8'h0E;
		16'h6BF1: out_word = 8'h00;
		16'h6BF2: out_word = 8'hCD;
		16'h6BF3: out_word = 8'h3A;
		16'h6BF4: out_word = 8'h2F;
		16'h6BF5: out_word = 8'hCD;
		16'h6BF6: out_word = 8'h34;
		16'h6BF7: out_word = 8'h2D;
		16'h6BF8: out_word = 8'h3A;
		16'h6BF9: out_word = 8'h02;
		16'h6BFA: out_word = 8'h41;
		16'h6BFB: out_word = 8'hCD;
		16'h6BFC: out_word = 8'hE5;
		16'h6BFD: out_word = 8'h2C;
		16'h6BFE: out_word = 8'h11;
		16'h6BFF: out_word = 8'h10;
		16'h6C00: out_word = 8'h41;
		16'h6C01: out_word = 8'h01;
		16'h6C02: out_word = 8'h10;
		16'h6C03: out_word = 8'h00;
		16'h6C04: out_word = 8'hEB;
		16'h6C05: out_word = 8'hED;
		16'h6C06: out_word = 8'hB0;
		16'h6C07: out_word = 8'hDB;
		16'h6C08: out_word = 8'h5F;
		16'h6C09: out_word = 8'h3D;
		16'h6C0A: out_word = 8'h5F;
		16'h6C0B: out_word = 8'h16;
		16'h6C0C: out_word = 8'h00;
		16'h6C0D: out_word = 8'h21;
		16'h6C0E: out_word = 8'h00;
		16'h6C0F: out_word = 8'h40;
		16'h6C10: out_word = 8'hCD;
		16'h6C11: out_word = 8'h73;
		16'h6C12: out_word = 8'h2D;
		16'h6C13: out_word = 8'h01;
		16'h6C14: out_word = 8'hFD;
		16'h6C15: out_word = 8'h7F;
		16'h6C16: out_word = 8'h3A;
		16'h6C17: out_word = 8'h01;
		16'h6C18: out_word = 8'h41;
		16'h6C19: out_word = 8'hED;
		16'h6C1A: out_word = 8'h79;
		16'h6C1B: out_word = 8'h2A;
		16'h6C1C: out_word = 8'h40;
		16'h6C1D: out_word = 8'h41;
		16'h6C1E: out_word = 8'hF9;
		16'h6C1F: out_word = 8'h21;
		16'h6C20: out_word = 8'h00;
		16'h6C21: out_word = 8'h40;
		16'h6C22: out_word = 8'h11;
		16'h6C23: out_word = 8'h0A;
		16'h6C24: out_word = 8'h00;
		16'h6C25: out_word = 8'hCD;
		16'h6C26: out_word = 8'h1B;
		16'h6C27: out_word = 8'h2F;
		16'h6C28: out_word = 8'h21;
		16'h6C29: out_word = 8'h00;
		16'h6C2A: out_word = 8'h41;
		16'h6C2B: out_word = 8'h11;
		16'h6C2C: out_word = 8'h0B;
		16'h6C2D: out_word = 8'h00;
		16'h6C2E: out_word = 8'hCD;
		16'h6C2F: out_word = 8'h1B;
		16'h6C30: out_word = 8'h2F;
		16'h6C31: out_word = 8'h3E;
		16'h6C32: out_word = 8'h3C;
		16'h6C33: out_word = 8'hF5;
		16'h6C34: out_word = 8'hC3;
		16'h6C35: out_word = 8'hBC;
		16'h6C36: out_word = 8'h2E;
		16'h6C37: out_word = 8'h78;
		16'h6C38: out_word = 8'h3D;
		16'h6C39: out_word = 8'h32;
		16'h6C3A: out_word = 8'h03;
		16'h6C3B: out_word = 8'h41;
		16'h6C3C: out_word = 8'h47;
		16'h6C3D: out_word = 8'h3A;
		16'h6C3E: out_word = 8'h01;
		16'h6C3F: out_word = 8'h41;
		16'h6C40: out_word = 8'hE6;
		16'h6C41: out_word = 8'h07;
		16'h6C42: out_word = 8'hB8;
		16'h6C43: out_word = 8'hC8;
		16'h6C44: out_word = 8'h3E;
		16'h6C45: out_word = 8'h02;
		16'h6C46: out_word = 8'hB8;
		16'h6C47: out_word = 8'hC8;
		16'h6C48: out_word = 8'h3A;
		16'h6C49: out_word = 8'h01;
		16'h6C4A: out_word = 8'h41;
		16'h6C4B: out_word = 8'hE6;
		16'h6C4C: out_word = 8'h08;
		16'h6C4D: out_word = 8'h28;
		16'h6C4E: out_word = 8'h06;
		16'h6C4F: out_word = 8'h78;
		16'h6C50: out_word = 8'hFE;
		16'h6C51: out_word = 8'h07;
		16'h6C52: out_word = 8'hC8;
		16'h6C53: out_word = 8'h18;
		16'h6C54: out_word = 8'h04;
		16'h6C55: out_word = 8'h78;
		16'h6C56: out_word = 8'hFE;
		16'h6C57: out_word = 8'h05;
		16'h6C58: out_word = 8'hC8;
		16'h6C59: out_word = 8'hCD;
		16'h6C5A: out_word = 8'h5D;
		16'h6C5B: out_word = 8'h2C;
		16'h6C5C: out_word = 8'hC9;
		16'h6C5D: out_word = 8'h21;
		16'h6C5E: out_word = 8'h01;
		16'h6C5F: out_word = 8'h41;
		16'h6C60: out_word = 8'h7E;
		16'h6C61: out_word = 8'hE6;
		16'h6C62: out_word = 8'hF8;
		16'h6C63: out_word = 8'h4F;
		16'h6C64: out_word = 8'h78;
		16'h6C65: out_word = 8'hB1;
		16'h6C66: out_word = 8'hC5;
		16'h6C67: out_word = 8'h01;
		16'h6C68: out_word = 8'hFD;
		16'h6C69: out_word = 8'h7F;
		16'h6C6A: out_word = 8'hED;
		16'h6C6B: out_word = 8'h79;
		16'h6C6C: out_word = 8'hC1;
		16'h6C6D: out_word = 8'h21;
		16'h6C6E: out_word = 8'h00;
		16'h6C6F: out_word = 8'hC0;
		16'h6C70: out_word = 8'h7E;
		16'h6C71: out_word = 8'hB7;
		16'h6C72: out_word = 8'h20;
		16'h6C73: out_word = 8'h06;
		16'h6C74: out_word = 8'h23;
		16'h6C75: out_word = 8'h7C;
		16'h6C76: out_word = 8'hB7;
		16'h6C77: out_word = 8'h20;
		16'h6C78: out_word = 8'hF7;
		16'h6C79: out_word = 8'hC9;
		16'h6C7A: out_word = 8'hCD;
		16'h6C7B: out_word = 8'h7E;
		16'h6C7C: out_word = 8'h2C;
		16'h6C7D: out_word = 8'hC9;
		16'h6C7E: out_word = 8'h0E;
		16'h6C7F: out_word = 8'h00;
		16'h6C80: out_word = 8'hCD;
		16'h6C81: out_word = 8'h3A;
		16'h6C82: out_word = 8'h2F;
		16'h6C83: out_word = 8'hCD;
		16'h6C84: out_word = 8'h2A;
		16'h6C85: out_word = 8'h2D;
		16'h6C86: out_word = 8'h3A;
		16'h6C87: out_word = 8'hE4;
		16'h6C88: out_word = 8'h40;
		16'h6C89: out_word = 8'h32;
		16'h6C8A: out_word = 8'h02;
		16'h6C8B: out_word = 8'h41;
		16'h6C8C: out_word = 8'h3C;
		16'h6C8D: out_word = 8'h32;
		16'h6C8E: out_word = 8'hE4;
		16'h6C8F: out_word = 8'h40;
		16'h6C90: out_word = 8'h2A;
		16'h6C91: out_word = 8'hE5;
		16'h6C92: out_word = 8'h40;
		16'h6C93: out_word = 8'h11;
		16'h6C94: out_word = 8'h40;
		16'h6C95: out_word = 8'h00;
		16'h6C96: out_word = 8'hED;
		16'h6C97: out_word = 8'h52;
		16'h6C98: out_word = 8'h22;
		16'h6C99: out_word = 8'hE5;
		16'h6C9A: out_word = 8'h40;
		16'h6C9B: out_word = 8'hD8;
		16'h6C9C: out_word = 8'h2A;
		16'h6C9D: out_word = 8'hE1;
		16'h6C9E: out_word = 8'h40;
		16'h6C9F: out_word = 8'h22;
		16'h6CA0: out_word = 8'h1E;
		16'h6CA1: out_word = 8'h41;
		16'h6CA2: out_word = 8'hCD;
		16'h6CA3: out_word = 8'h1E;
		16'h6CA4: out_word = 8'h2D;
		16'h6CA5: out_word = 8'h3E;
		16'h6CA6: out_word = 8'h40;
		16'h6CA7: out_word = 8'h32;
		16'h6CA8: out_word = 8'h1D;
		16'h6CA9: out_word = 8'h41;
		16'h6CAA: out_word = 8'h21;
		16'h6CAB: out_word = 8'h00;
		16'h6CAC: out_word = 8'hC0;
		16'h6CAD: out_word = 8'h22;
		16'h6CAE: out_word = 8'h19;
		16'h6CAF: out_word = 8'h41;
		16'h6CB0: out_word = 8'h21;
		16'h6CB1: out_word = 8'h00;
		16'h6CB2: out_word = 8'h40;
		16'h6CB3: out_word = 8'h22;
		16'h6CB4: out_word = 8'h1B;
		16'h6CB5: out_word = 8'h41;
		16'h6CB6: out_word = 8'hED;
		16'h6CB7: out_word = 8'h5B;
		16'h6CB8: out_word = 8'hE1;
		16'h6CB9: out_word = 8'h40;
		16'h6CBA: out_word = 8'hCD;
		16'h6CBB: out_word = 8'h3E;
		16'h6CBC: out_word = 8'h2D;
		16'h6CBD: out_word = 8'hED;
		16'h6CBE: out_word = 8'h53;
		16'h6CBF: out_word = 8'hE1;
		16'h6CC0: out_word = 8'h40;
		16'h6CC1: out_word = 8'h0E;
		16'h6CC2: out_word = 8'h00;
		16'h6CC3: out_word = 8'hCD;
		16'h6CC4: out_word = 8'h3A;
		16'h6CC5: out_word = 8'h2F;
		16'h6CC6: out_word = 8'hCD;
		16'h6CC7: out_word = 8'h34;
		16'h6CC8: out_word = 8'h2D;
		16'h6CC9: out_word = 8'h3A;
		16'h6CCA: out_word = 8'h02;
		16'h6CCB: out_word = 8'h41;
		16'h6CCC: out_word = 8'hCD;
		16'h6CCD: out_word = 8'hE5;
		16'h6CCE: out_word = 8'h2C;
		16'h6CCF: out_word = 8'h11;
		16'h6CD0: out_word = 8'h10;
		16'h6CD1: out_word = 8'h41;
		16'h6CD2: out_word = 8'h01;
		16'h6CD3: out_word = 8'h10;
		16'h6CD4: out_word = 8'h00;
		16'h6CD5: out_word = 8'hEB;
		16'h6CD6: out_word = 8'hED;
		16'h6CD7: out_word = 8'hB0;
		16'h6CD8: out_word = 8'hDB;
		16'h6CD9: out_word = 8'h5F;
		16'h6CDA: out_word = 8'h3D;
		16'h6CDB: out_word = 8'h5F;
		16'h6CDC: out_word = 8'h16;
		16'h6CDD: out_word = 8'h00;
		16'h6CDE: out_word = 8'h21;
		16'h6CDF: out_word = 8'h00;
		16'h6CE0: out_word = 8'h40;
		16'h6CE1: out_word = 8'hCD;
		16'h6CE2: out_word = 8'h73;
		16'h6CE3: out_word = 8'h2D;
		16'h6CE4: out_word = 8'hC9;
		16'h6CE5: out_word = 8'h4F;
		16'h6CE6: out_word = 8'hE6;
		16'h6CE7: out_word = 8'hF0;
		16'h6CE8: out_word = 8'h0F;
		16'h6CE9: out_word = 8'h0F;
		16'h6CEA: out_word = 8'h0F;
		16'h6CEB: out_word = 8'h0F;
		16'h6CEC: out_word = 8'h47;
		16'h6CED: out_word = 8'hC5;
		16'h6CEE: out_word = 8'h58;
		16'h6CEF: out_word = 8'h16;
		16'h6CF0: out_word = 8'h00;
		16'h6CF1: out_word = 8'h21;
		16'h6CF2: out_word = 8'h00;
		16'h6CF3: out_word = 8'h40;
		16'h6CF4: out_word = 8'hD5;
		16'h6CF5: out_word = 8'hCD;
		16'h6CF6: out_word = 8'h1B;
		16'h6CF7: out_word = 8'h2F;
		16'h6CF8: out_word = 8'hD1;
		16'h6CF9: out_word = 8'hC1;
		16'h6CFA: out_word = 8'h06;
		16'h6CFB: out_word = 8'h00;
		16'h6CFC: out_word = 8'h79;
		16'h6CFD: out_word = 8'hE6;
		16'h6CFE: out_word = 8'h0F;
		16'h6CFF: out_word = 8'h07;
		16'h6D00: out_word = 8'h07;
		16'h6D01: out_word = 8'h07;
		16'h6D02: out_word = 8'h07;
		16'h6D03: out_word = 8'h21;
		16'h6D04: out_word = 8'h00;
		16'h6D05: out_word = 8'h40;
		16'h6D06: out_word = 8'h85;
		16'h6D07: out_word = 8'h6F;
		16'h6D08: out_word = 8'hC9;
		16'h6D09: out_word = 8'h21;
		16'h6D0A: out_word = 8'h10;
		16'h6D0B: out_word = 8'h41;
		16'h6D0C: out_word = 8'h06;
		16'h6D0D: out_word = 8'h09;
		16'h6D0E: out_word = 8'h36;
		16'h6D0F: out_word = 8'h20;
		16'h6D10: out_word = 8'h23;
		16'h6D11: out_word = 8'h10;
		16'h6D12: out_word = 8'hFB;
		16'h6D13: out_word = 8'h3E;
		16'h6D14: out_word = 8'h40;
		16'h6D15: out_word = 8'h32;
		16'h6D16: out_word = 8'h10;
		16'h6D17: out_word = 8'h41;
		16'h6D18: out_word = 8'h3E;
		16'h6D19: out_word = 8'h43;
		16'h6D1A: out_word = 8'h32;
		16'h6D1B: out_word = 8'h18;
		16'h6D1C: out_word = 8'h41;
		16'h6D1D: out_word = 8'hC9;
		16'h6D1E: out_word = 8'hCD;
		16'h6D1F: out_word = 8'h09;
		16'h6D20: out_word = 8'h2D;
		16'h6D21: out_word = 8'h3A;
		16'h6D22: out_word = 8'h03;
		16'h6D23: out_word = 8'h41;
		16'h6D24: out_word = 8'hC6;
		16'h6D25: out_word = 8'h30;
		16'h6D26: out_word = 8'h32;
		16'h6D27: out_word = 8'h11;
		16'h6D28: out_word = 8'h41;
		16'h6D29: out_word = 8'hC9;
		16'h6D2A: out_word = 8'h21;
		16'h6D2B: out_word = 8'h00;
		16'h6D2C: out_word = 8'h40;
		16'h6D2D: out_word = 8'h11;
		16'h6D2E: out_word = 8'h08;
		16'h6D2F: out_word = 8'h00;
		16'h6D30: out_word = 8'hCD;
		16'h6D31: out_word = 8'h1B;
		16'h6D32: out_word = 8'h2F;
		16'h6D33: out_word = 8'hC9;
		16'h6D34: out_word = 8'h21;
		16'h6D35: out_word = 8'h00;
		16'h6D36: out_word = 8'h40;
		16'h6D37: out_word = 8'h11;
		16'h6D38: out_word = 8'h08;
		16'h6D39: out_word = 8'h00;
		16'h6D3A: out_word = 8'hCD;
		16'h6D3B: out_word = 8'h73;
		16'h6D3C: out_word = 8'h2D;
		16'h6D3D: out_word = 8'hC9;
		16'h6D3E: out_word = 8'hCD;
		16'h6D3F: out_word = 8'h65;
		16'h6D40: out_word = 8'h2F;
		16'h6D41: out_word = 8'h4A;
		16'h6D42: out_word = 8'hCD;
		16'h6D43: out_word = 8'h3A;
		16'h6D44: out_word = 8'h2F;
		16'h6D45: out_word = 8'h21;
		16'h6D46: out_word = 8'h00;
		16'h6D47: out_word = 8'hC0;
		16'h6D48: out_word = 8'h06;
		16'h6D49: out_word = 8'h40;
		16'h6D4A: out_word = 8'h18;
		16'h6D4B: out_word = 8'h0C;
		16'h6D4C: out_word = 8'hCD;
		16'h6D4D: out_word = 8'h65;
		16'h6D4E: out_word = 8'h2F;
		16'h6D4F: out_word = 8'h4A;
		16'h6D50: out_word = 8'hCD;
		16'h6D51: out_word = 8'h3A;
		16'h6D52: out_word = 8'h2F;
		16'h6D53: out_word = 8'h21;
		16'h6D54: out_word = 8'h00;
		16'h6D55: out_word = 8'h40;
		16'h6D56: out_word = 8'h06;
		16'h6D57: out_word = 8'hC0;
		16'h6D58: out_word = 8'hC5;
		16'h6D59: out_word = 8'hD5;
		16'h6D5A: out_word = 8'hCD;
		16'h6D5B: out_word = 8'h73;
		16'h6D5C: out_word = 8'h2D;
		16'h6D5D: out_word = 8'h11;
		16'h6D5E: out_word = 8'h00;
		16'h6D5F: out_word = 8'h01;
		16'h6D60: out_word = 8'h19;
		16'h6D61: out_word = 8'hD1;
		16'h6D62: out_word = 8'h1C;
		16'h6D63: out_word = 8'h7B;
		16'h6D64: out_word = 8'hFE;
		16'h6D65: out_word = 8'h10;
		16'h6D66: out_word = 8'h20;
		16'h6D67: out_word = 8'h07;
		16'h6D68: out_word = 8'h1E;
		16'h6D69: out_word = 8'h00;
		16'h6D6A: out_word = 8'h14;
		16'h6D6B: out_word = 8'h4A;
		16'h6D6C: out_word = 8'hCD;
		16'h6D6D: out_word = 8'h3A;
		16'h6D6E: out_word = 8'h2F;
		16'h6D6F: out_word = 8'hC1;
		16'h6D70: out_word = 8'h10;
		16'h6D71: out_word = 8'hE6;
		16'h6D72: out_word = 8'hC9;
		16'h6D73: out_word = 8'h7B;
		16'h6D74: out_word = 8'h3C;
		16'h6D75: out_word = 8'hD3;
		16'h6D76: out_word = 8'h5F;
		16'h6D77: out_word = 8'hE5;
		16'h6D78: out_word = 8'h16;
		16'h6D79: out_word = 8'h14;
		16'h6D7A: out_word = 8'hD5;
		16'h6D7B: out_word = 8'hF3;
		16'h6D7C: out_word = 8'h0E;
		16'h6D7D: out_word = 8'h7F;
		16'h6D7E: out_word = 8'h3E;
		16'h6D7F: out_word = 8'hA0;
		16'h6D80: out_word = 8'hD3;
		16'h6D81: out_word = 8'h1F;
		16'h6D82: out_word = 8'hCD;
		16'h6D83: out_word = 8'hCA;
		16'h6D84: out_word = 8'h3F;
		16'h6D85: out_word = 8'hD1;
		16'h6D86: out_word = 8'hE1;
		16'h6D87: out_word = 8'hDB;
		16'h6D88: out_word = 8'h1F;
		16'h6D89: out_word = 8'hE6;
		16'h6D8A: out_word = 8'h7F;
		16'h6D8B: out_word = 8'hC8;
		16'h6D8C: out_word = 8'h15;
		16'h6D8D: out_word = 8'hE5;
		16'h6D8E: out_word = 8'hD5;
		16'h6D8F: out_word = 8'h20;
		16'h6D90: out_word = 8'hEA;
		16'h6D91: out_word = 8'h76;
		16'h6D92: out_word = 8'h2A;
		16'h6D93: out_word = 8'hE6;
		16'h6D94: out_word = 8'h5C;
		16'h6D95: out_word = 8'hED;
		16'h6D96: out_word = 8'h5B;
		16'h6D97: out_word = 8'hEB;
		16'h6D98: out_word = 8'h5C;
		16'h6D99: out_word = 8'h3A;
		16'h6D9A: out_word = 8'hEA;
		16'h6D9B: out_word = 8'h5C;
		16'h6D9C: out_word = 8'h47;
		16'h6D9D: out_word = 8'hCD;
		16'h6D9E: out_word = 8'h3D;
		16'h6D9F: out_word = 8'h1E;
		16'h6DA0: out_word = 8'hC9;
		16'h6DA1: out_word = 8'hCD;
		16'h6DA2: out_word = 8'hDF;
		16'h6DA3: out_word = 8'h1D;
		16'h6DA4: out_word = 8'hCD;
		16'h6DA5: out_word = 8'h75;
		16'h6DA6: out_word = 8'h1D;
		16'h6DA7: out_word = 8'hCD;
		16'h6DA8: out_word = 8'h2E;
		16'h6DA9: out_word = 8'h10;
		16'h6DAA: out_word = 8'hCD;
		16'h6DAB: out_word = 8'h57;
		16'h6DAC: out_word = 8'h1C;
		16'h6DAD: out_word = 8'hED;
		16'h6DAE: out_word = 8'h43;
		16'h6DAF: out_word = 8'h20;
		16'h6DB0: out_word = 8'h40;
		16'h6DB1: out_word = 8'h79;
		16'h6DB2: out_word = 8'hFE;
		16'h6DB3: out_word = 8'h08;
		16'h6DB4: out_word = 8'h30;
		16'h6DB5: out_word = 8'h1C;
		16'h6DB6: out_word = 8'hCD;
		16'h6DB7: out_word = 8'h05;
		16'h6DB8: out_word = 8'h04;
		16'h6DB9: out_word = 8'hCD;
		16'h6DBA: out_word = 8'hB3;
		16'h6DBB: out_word = 8'h1C;
		16'h6DBC: out_word = 8'hC2;
		16'h6DBD: out_word = 8'hD9;
		16'h6DBE: out_word = 8'h03;
		16'h6DBF: out_word = 8'h21;
		16'h6DC0: out_word = 8'hDD;
		16'h6DC1: out_word = 8'h5C;
		16'h6DC2: out_word = 8'hED;
		16'h6DC3: out_word = 8'h4B;
		16'h6DC4: out_word = 8'h20;
		16'h6DC5: out_word = 8'h40;
		16'h6DC6: out_word = 8'h09;
		16'h6DC7: out_word = 8'h36;
		16'h6DC8: out_word = 8'h38;
		16'h6DC9: out_word = 8'hE5;
		16'h6DCA: out_word = 8'hCD;
		16'h6DCB: out_word = 8'hB3;
		16'h6DCC: out_word = 8'h1C;
		16'h6DCD: out_word = 8'hE1;
		16'h6DCE: out_word = 8'h28;
		16'h6DCF: out_word = 8'h08;
		16'h6DD0: out_word = 8'h36;
		16'h6DD1: out_word = 8'h20;
		16'h6DD2: out_word = 8'hCD;
		16'h6DD3: out_word = 8'hB3;
		16'h6DD4: out_word = 8'h1C;
		16'h6DD5: out_word = 8'hC3;
		16'h6DD6: out_word = 8'h33;
		16'h6DD7: out_word = 8'h2E;
		16'h6DD8: out_word = 8'hCD;
		16'h6DD9: out_word = 8'h5D;
		16'h6DDA: out_word = 8'h16;
		16'h6DDB: out_word = 8'hCD;
		16'h6DDC: out_word = 8'h92;
		16'h6DDD: out_word = 8'h2D;
		16'h6DDE: out_word = 8'h31;
		16'h6DDF: out_word = 8'hFF;
		16'h6DE0: out_word = 8'h40;
		16'h6DE1: out_word = 8'h06;
		16'h6DE2: out_word = 8'h08;
		16'h6DE3: out_word = 8'hC5;
		16'h6DE4: out_word = 8'h78;
		16'h6DE5: out_word = 8'h01;
		16'h6DE6: out_word = 8'hFD;
		16'h6DE7: out_word = 8'h7F;
		16'h6DE8: out_word = 8'h3D;
		16'h6DE9: out_word = 8'hF5;
		16'h6DEA: out_word = 8'hF6;
		16'h6DEB: out_word = 8'h10;
		16'h6DEC: out_word = 8'hED;
		16'h6DED: out_word = 8'h79;
		16'h6DEE: out_word = 8'hF1;
		16'h6DEF: out_word = 8'hC6;
		16'h6DF0: out_word = 8'h30;
		16'h6DF1: out_word = 8'h21;
		16'h6DF2: out_word = 8'hDD;
		16'h6DF3: out_word = 8'h5C;
		16'h6DF4: out_word = 8'hED;
		16'h6DF5: out_word = 8'h4B;
		16'h6DF6: out_word = 8'h20;
		16'h6DF7: out_word = 8'h40;
		16'h6DF8: out_word = 8'h09;
		16'h6DF9: out_word = 8'h77;
		16'h6DFA: out_word = 8'hCD;
		16'h6DFB: out_word = 8'hB3;
		16'h6DFC: out_word = 8'h1C;
		16'h6DFD: out_word = 8'h20;
		16'h6DFE: out_word = 8'h06;
		16'h6DFF: out_word = 8'hCD;
		16'h6E00: out_word = 8'h5D;
		16'h6E01: out_word = 8'h16;
		16'h6E02: out_word = 8'hCD;
		16'h6E03: out_word = 8'h92;
		16'h6E04: out_word = 8'h2D;
		16'h6E05: out_word = 8'hC1;
		16'h6E06: out_word = 8'h10;
		16'h6E07: out_word = 8'hDB;
		16'h6E08: out_word = 8'h3E;
		16'h6E09: out_word = 8'h20;
		16'h6E0A: out_word = 8'h21;
		16'h6E0B: out_word = 8'hDD;
		16'h6E0C: out_word = 8'h5C;
		16'h6E0D: out_word = 8'hED;
		16'h6E0E: out_word = 8'h4B;
		16'h6E0F: out_word = 8'h20;
		16'h6E10: out_word = 8'h40;
		16'h6E11: out_word = 8'h09;
		16'h6E12: out_word = 8'h77;
		16'h6E13: out_word = 8'hCD;
		16'h6E14: out_word = 8'hB3;
		16'h6E15: out_word = 8'h1C;
		16'h6E16: out_word = 8'hCD;
		16'h6E17: out_word = 8'h5D;
		16'h6E18: out_word = 8'h16;
		16'h6E19: out_word = 8'hC5;
		16'h6E1A: out_word = 8'hF5;
		16'h6E1B: out_word = 8'h01;
		16'h6E1C: out_word = 8'hFD;
		16'h6E1D: out_word = 8'h7F;
		16'h6E1E: out_word = 8'h3A;
		16'h6E1F: out_word = 8'h01;
		16'h6E20: out_word = 8'h41;
		16'h6E21: out_word = 8'hED;
		16'h6E22: out_word = 8'h79;
		16'h6E23: out_word = 8'hF1;
		16'h6E24: out_word = 8'hC1;
		16'h6E25: out_word = 8'h18;
		16'h6E26: out_word = 8'h12;
		16'h6E27: out_word = 8'hCD;
		16'h6E28: out_word = 8'hDF;
		16'h6E29: out_word = 8'h1D;
		16'h6E2A: out_word = 8'hCD;
		16'h6E2B: out_word = 8'h75;
		16'h6E2C: out_word = 8'h1D;
		16'h6E2D: out_word = 8'hCD;
		16'h6E2E: out_word = 8'h2E;
		16'h6E2F: out_word = 8'h10;
		16'h6E30: out_word = 8'hCD;
		16'h6E31: out_word = 8'h2F;
		16'h6E32: out_word = 8'h29;
		16'h6E33: out_word = 8'hC2;
		16'h6E34: out_word = 8'hD9;
		16'h6E35: out_word = 8'h03;
		16'h6E36: out_word = 8'hCD;
		16'h6E37: out_word = 8'h5D;
		16'h6E38: out_word = 8'h16;
		16'h6E39: out_word = 8'h3A;
		16'h6E3A: out_word = 8'hDD;
		16'h6E3B: out_word = 8'h5C;
		16'h6E3C: out_word = 8'hFE;
		16'h6E3D: out_word = 8'h24;
		16'h6E3E: out_word = 8'hF3;
		16'h6E3F: out_word = 8'h20;
		16'h6E40: out_word = 8'h02;
		16'h6E41: out_word = 8'hED;
		16'h6E42: out_word = 8'h5E;
		16'h6E43: out_word = 8'h31;
		16'h6E44: out_word = 8'hF0;
		16'h6E45: out_word = 8'h40;
		16'h6E46: out_word = 8'hCD;
		16'h6E47: out_word = 8'h11;
		16'h6E48: out_word = 8'h3E;
		16'h6E49: out_word = 8'h32;
		16'h6E4A: out_word = 8'h10;
		16'h6E4B: out_word = 8'h40;
		16'h6E4C: out_word = 8'h3A;
		16'h6E4D: out_word = 8'h16;
		16'h6E4E: out_word = 8'h5D;
		16'h6E4F: out_word = 8'h32;
		16'h6E50: out_word = 8'h11;
		16'h6E51: out_word = 8'h40;
		16'h6E52: out_word = 8'h2A;
		16'h6E53: out_word = 8'hE6;
		16'h6E54: out_word = 8'h5C;
		16'h6E55: out_word = 8'hE5;
		16'h6E56: out_word = 8'hED;
		16'h6E57: out_word = 8'h5B;
		16'h6E58: out_word = 8'hEB;
		16'h6E59: out_word = 8'h5C;
		16'h6E5A: out_word = 8'hD5;
		16'h6E5B: out_word = 8'h1C;
		16'h6E5C: out_word = 8'h7B;
		16'h6E5D: out_word = 8'hFE;
		16'h6E5E: out_word = 8'h10;
		16'h6E5F: out_word = 8'h20;
		16'h6E60: out_word = 8'h03;
		16'h6E61: out_word = 8'h1E;
		16'h6E62: out_word = 8'h00;
		16'h6E63: out_word = 8'h14;
		16'h6E64: out_word = 8'h4A;
		16'h6E65: out_word = 8'hCD;
		16'h6E66: out_word = 8'h07;
		16'h6E67: out_word = 8'h2F;
		16'h6E68: out_word = 8'h3A;
		16'h6E69: out_word = 8'h10;
		16'h6E6A: out_word = 8'h40;
		16'h6E6B: out_word = 8'hE6;
		16'h6E6C: out_word = 8'h02;
		16'h6E6D: out_word = 8'hC4;
		16'h6E6E: out_word = 8'h0F;
		16'h6E6F: out_word = 8'h2F;
		16'h6E70: out_word = 8'h79;
		16'h6E71: out_word = 8'hCD;
		16'h6E72: out_word = 8'h50;
		16'h6E73: out_word = 8'h2F;
		16'h6E74: out_word = 8'h21;
		16'h6E75: out_word = 8'h00;
		16'h6E76: out_word = 8'h41;
		16'h6E77: out_word = 8'h06;
		16'h6E78: out_word = 8'hBF;
		16'h6E79: out_word = 8'hC5;
		16'h6E7A: out_word = 8'hD5;
		16'h6E7B: out_word = 8'hCD;
		16'h6E7C: out_word = 8'h1B;
		16'h6E7D: out_word = 8'h2F;
		16'h6E7E: out_word = 8'h11;
		16'h6E7F: out_word = 8'h00;
		16'h6E80: out_word = 8'h01;
		16'h6E81: out_word = 8'h19;
		16'h6E82: out_word = 8'hD1;
		16'h6E83: out_word = 8'h1C;
		16'h6E84: out_word = 8'h7B;
		16'h6E85: out_word = 8'hFE;
		16'h6E86: out_word = 8'h10;
		16'h6E87: out_word = 8'h20;
		16'h6E88: out_word = 8'h13;
		16'h6E89: out_word = 8'h1E;
		16'h6E8A: out_word = 8'h00;
		16'h6E8B: out_word = 8'h14;
		16'h6E8C: out_word = 8'h4A;
		16'h6E8D: out_word = 8'hCD;
		16'h6E8E: out_word = 8'h07;
		16'h6E8F: out_word = 8'h2F;
		16'h6E90: out_word = 8'h3A;
		16'h6E91: out_word = 8'h10;
		16'h6E92: out_word = 8'h40;
		16'h6E93: out_word = 8'hE6;
		16'h6E94: out_word = 8'h02;
		16'h6E95: out_word = 8'hC4;
		16'h6E96: out_word = 8'h0F;
		16'h6E97: out_word = 8'h2F;
		16'h6E98: out_word = 8'h79;
		16'h6E99: out_word = 8'hCD;
		16'h6E9A: out_word = 8'h50;
		16'h6E9B: out_word = 8'h2F;
		16'h6E9C: out_word = 8'hC1;
		16'h6E9D: out_word = 8'h10;
		16'h6E9E: out_word = 8'hDA;
		16'h6E9F: out_word = 8'hD1;
		16'h6EA0: out_word = 8'hE1;
		16'h6EA1: out_word = 8'hF9;
		16'h6EA2: out_word = 8'h3A;
		16'h6EA3: out_word = 8'h11;
		16'h6EA4: out_word = 8'h40;
		16'h6EA5: out_word = 8'hF5;
		16'h6EA6: out_word = 8'h4A;
		16'h6EA7: out_word = 8'hCD;
		16'h6EA8: out_word = 8'h07;
		16'h6EA9: out_word = 8'h2F;
		16'h6EAA: out_word = 8'h3A;
		16'h6EAB: out_word = 8'h10;
		16'h6EAC: out_word = 8'h40;
		16'h6EAD: out_word = 8'hE6;
		16'h6EAE: out_word = 8'h02;
		16'h6EAF: out_word = 8'hC4;
		16'h6EB0: out_word = 8'h0F;
		16'h6EB1: out_word = 8'h2F;
		16'h6EB2: out_word = 8'h79;
		16'h6EB3: out_word = 8'hCD;
		16'h6EB4: out_word = 8'h50;
		16'h6EB5: out_word = 8'h2F;
		16'h6EB6: out_word = 8'h21;
		16'h6EB7: out_word = 8'h00;
		16'h6EB8: out_word = 8'h40;
		16'h6EB9: out_word = 8'hCD;
		16'h6EBA: out_word = 8'h1B;
		16'h6EBB: out_word = 8'h2F;
		16'h6EBC: out_word = 8'hF1;
		16'h6EBD: out_word = 8'h08;
		16'h6EBE: out_word = 8'hF1;
		16'h6EBF: out_word = 8'hC3;
		16'h6EC0: out_word = 8'h0A;
		16'h6EC1: out_word = 8'h0A;
		16'h6EC2: out_word = 8'hED;
		16'h6EC3: out_word = 8'h47;
		16'h6EC4: out_word = 8'hF3;
		16'h6EC5: out_word = 8'h3E;
		16'h6EC6: out_word = 8'hFF;
		16'h6EC7: out_word = 8'hE2;
		16'h6EC8: out_word = 8'hCC;
		16'h6EC9: out_word = 8'h2E;
		16'h6ECA: out_word = 8'h3E;
		16'h6ECB: out_word = 8'h00;
		16'h6ECC: out_word = 8'h32;
		16'h6ECD: out_word = 8'h00;
		16'h6ECE: out_word = 8'h5C;
		16'h6ECF: out_word = 8'hF1;
		16'h6ED0: out_word = 8'hE1;
		16'h6ED1: out_word = 8'hD1;
		16'h6ED2: out_word = 8'hC1;
		16'h6ED3: out_word = 8'hD9;
		16'h6ED4: out_word = 8'h08;
		16'h6ED5: out_word = 8'hFD;
		16'h6ED6: out_word = 8'hE1;
		16'h6ED7: out_word = 8'hDD;
		16'h6ED8: out_word = 8'hE1;
		16'h6ED9: out_word = 8'hE1;
		16'h6EDA: out_word = 8'hD1;
		16'h6EDB: out_word = 8'hC1;
		16'h6EDC: out_word = 8'h3A;
		16'h6EDD: out_word = 8'h48;
		16'h6EDE: out_word = 8'h5C;
		16'h6EDF: out_word = 8'hE6;
		16'h6EE0: out_word = 8'h38;
		16'h6EE1: out_word = 8'h0F;
		16'h6EE2: out_word = 8'h0F;
		16'h6EE3: out_word = 8'h0F;
		16'h6EE4: out_word = 8'hD3;
		16'h6EE5: out_word = 8'hFE;
		16'h6EE6: out_word = 8'h3A;
		16'h6EE7: out_word = 8'h08;
		16'h6EE8: out_word = 8'h5B;
		16'h6EE9: out_word = 8'hFE;
		16'h6EEA: out_word = 8'hEE;
		16'h6EEB: out_word = 8'h20;
		16'h6EEC: out_word = 8'h0A;
		16'h6EED: out_word = 8'hC5;
		16'h6EEE: out_word = 8'h01;
		16'h6EEF: out_word = 8'hFD;
		16'h6EF0: out_word = 8'h7F;
		16'h6EF1: out_word = 8'h3A;
		16'h6EF2: out_word = 8'h5C;
		16'h6EF3: out_word = 8'h5B;
		16'h6EF4: out_word = 8'hED;
		16'h6EF5: out_word = 8'h79;
		16'h6EF6: out_word = 8'hC1;
		16'h6EF7: out_word = 8'h3A;
		16'h6EF8: out_word = 8'h00;
		16'h6EF9: out_word = 8'h5C;
		16'h6EFA: out_word = 8'hB7;
		16'h6EFB: out_word = 8'h3E;
		16'h6EFC: out_word = 8'hC9;
		16'h6EFD: out_word = 8'h32;
		16'h6EFE: out_word = 8'h00;
		16'h6EFF: out_word = 8'h5C;
		16'h6F00: out_word = 8'h20;
		16'h6F01: out_word = 8'h01;
		16'h6F02: out_word = 8'hFB;
		16'h6F03: out_word = 8'hC3;
		16'h6F04: out_word = 8'h11;
		16'h6F05: out_word = 8'h0A;
		16'h6F06: out_word = 8'h00;
		16'h6F07: out_word = 8'h3A;
		16'h6F08: out_word = 8'h11;
		16'h6F09: out_word = 8'h40;
		16'h6F0A: out_word = 8'hF6;
		16'h6F0B: out_word = 8'h3C;
		16'h6F0C: out_word = 8'hD3;
		16'h6F0D: out_word = 8'hFF;
		16'h6F0E: out_word = 8'hC9;
		16'h6F0F: out_word = 8'h79;
		16'h6F10: out_word = 8'hB7;
		16'h6F11: out_word = 8'h1F;
		16'h6F12: out_word = 8'h4F;
		16'h6F13: out_word = 8'hD0;
		16'h6F14: out_word = 8'h3A;
		16'h6F15: out_word = 8'h11;
		16'h6F16: out_word = 8'h40;
		16'h6F17: out_word = 8'hE6;
		16'h6F18: out_word = 8'h6F;
		16'h6F19: out_word = 8'h18;
		16'h6F1A: out_word = 8'hF1;
		16'h6F1B: out_word = 8'h7B;
		16'h6F1C: out_word = 8'h3C;
		16'h6F1D: out_word = 8'hD3;
		16'h6F1E: out_word = 8'h5F;
		16'h6F1F: out_word = 8'hE5;
		16'h6F20: out_word = 8'h16;
		16'h6F21: out_word = 8'h14;
		16'h6F22: out_word = 8'hD5;
		16'h6F23: out_word = 8'hF3;
		16'h6F24: out_word = 8'h0E;
		16'h6F25: out_word = 8'h7F;
		16'h6F26: out_word = 8'h3E;
		16'h6F27: out_word = 8'h80;
		16'h6F28: out_word = 8'hD3;
		16'h6F29: out_word = 8'h1F;
		16'h6F2A: out_word = 8'hCD;
		16'h6F2B: out_word = 8'hE5;
		16'h6F2C: out_word = 8'h3F;
		16'h6F2D: out_word = 8'hD1;
		16'h6F2E: out_word = 8'hE1;
		16'h6F2F: out_word = 8'hDB;
		16'h6F30: out_word = 8'h1F;
		16'h6F31: out_word = 8'hE6;
		16'h6F32: out_word = 8'h7F;
		16'h6F33: out_word = 8'hC8;
		16'h6F34: out_word = 8'h15;
		16'h6F35: out_word = 8'hE5;
		16'h6F36: out_word = 8'hD5;
		16'h6F37: out_word = 8'h20;
		16'h6F38: out_word = 8'hEA;
		16'h6F39: out_word = 8'h76;
		16'h6F3A: out_word = 8'h3E;
		16'h6F3B: out_word = 8'h3C;
		16'h6F3C: out_word = 8'hD3;
		16'h6F3D: out_word = 8'hFF;
		16'h6F3E: out_word = 8'h3A;
		16'h6F3F: out_word = 8'h00;
		16'h6F40: out_word = 8'h5C;
		16'h6F41: out_word = 8'hE6;
		16'h6F42: out_word = 8'h08;
		16'h6F43: out_word = 8'h20;
		16'h6F44: out_word = 8'h0A;
		16'h6F45: out_word = 8'h79;
		16'h6F46: out_word = 8'hB7;
		16'h6F47: out_word = 8'h1F;
		16'h6F48: out_word = 8'h4F;
		16'h6F49: out_word = 8'h30;
		16'h6F4A: out_word = 8'h04;
		16'h6F4B: out_word = 8'h3E;
		16'h6F4C: out_word = 8'h2C;
		16'h6F4D: out_word = 8'hD3;
		16'h6F4E: out_word = 8'hFF;
		16'h6F4F: out_word = 8'h79;
		16'h6F50: out_word = 8'hD3;
		16'h6F51: out_word = 8'h7F;
		16'h6F52: out_word = 8'hCD;
		16'h6F53: out_word = 8'h30;
		16'h6F54: out_word = 8'h3D;
		16'h6F55: out_word = 8'h3E;
		16'h6F56: out_word = 8'h18;
		16'h6F57: out_word = 8'hD3;
		16'h6F58: out_word = 8'h1F;
		16'h6F59: out_word = 8'hDB;
		16'h6F5A: out_word = 8'hFF;
		16'h6F5B: out_word = 8'hE6;
		16'h6F5C: out_word = 8'h80;
		16'h6F5D: out_word = 8'h28;
		16'h6F5E: out_word = 8'hFA;
		16'h6F5F: out_word = 8'hC5;
		16'h6F60: out_word = 8'hCD;
		16'h6F61: out_word = 8'hFD;
		16'h6F62: out_word = 8'h3D;
		16'h6F63: out_word = 8'hC1;
		16'h6F64: out_word = 8'hC9;
		16'h6F65: out_word = 8'h3E;
		16'h6F66: out_word = 8'h08;
		16'h6F67: out_word = 8'h18;
		16'h6F68: out_word = 8'hEE;
		16'h6F69: out_word = 8'h2A;
		16'h6F6A: out_word = 8'h1C;
		16'h6F6B: out_word = 8'h5D;
		16'h6F6C: out_word = 8'h2B;
		16'h6F6D: out_word = 8'h2B;
		16'h6F6E: out_word = 8'hF9;
		16'h6F6F: out_word = 8'hC3;
		16'h6F70: out_word = 8'h2F;
		16'h6F71: out_word = 8'h1D;
		16'h6F72: out_word = 8'h22;
		16'h6F73: out_word = 8'h02;
		16'h6F74: out_word = 8'h5D;
		16'h6F75: out_word = 8'hED;
		16'h6F76: out_word = 8'h53;
		16'h6F77: out_word = 8'h04;
		16'h6F78: out_word = 8'h5D;
		16'h6F79: out_word = 8'hE1;
		16'h6F7A: out_word = 8'h5E;
		16'h6F7B: out_word = 8'h23;
		16'h6F7C: out_word = 8'h56;
		16'h6F7D: out_word = 8'h23;
		16'h6F7E: out_word = 8'hE5;
		16'h6F7F: out_word = 8'h21;
		16'h6F80: out_word = 8'h2F;
		16'h6F81: out_word = 8'h3D;
		16'h6F82: out_word = 8'hE5;
		16'h6F83: out_word = 8'hD5;
		16'h6F84: out_word = 8'h21;
		16'h6F85: out_word = 8'hC2;
		16'h6F86: out_word = 8'h5C;
		16'h6F87: out_word = 8'hE5;
		16'h6F88: out_word = 8'h2A;
		16'h6F89: out_word = 8'h02;
		16'h6F8A: out_word = 8'h5D;
		16'h6F8B: out_word = 8'hED;
		16'h6F8C: out_word = 8'h5B;
		16'h6F8D: out_word = 8'h04;
		16'h6F8E: out_word = 8'h5D;
		16'h6F8F: out_word = 8'hC9;
		16'h6F90: out_word = 8'h21;
		16'h6F91: out_word = 8'hFF;
		16'h6F92: out_word = 8'hFF;
		16'h6F93: out_word = 8'h22;
		16'h6F94: out_word = 8'hFA;
		16'h6F95: out_word = 8'h5C;
		16'h6F96: out_word = 8'h22;
		16'h6F97: out_word = 8'hFC;
		16'h6F98: out_word = 8'h5C;
		16'h6F99: out_word = 8'h22;
		16'h6F9A: out_word = 8'hC8;
		16'h6F9B: out_word = 8'h5C;
		16'h6F9C: out_word = 8'h22;
		16'h6F9D: out_word = 8'hCA;
		16'h6F9E: out_word = 8'h5C;
		16'h6F9F: out_word = 8'hAF;
		16'h6FA0: out_word = 8'h32;
		16'h6FA1: out_word = 8'h17;
		16'h6FA2: out_word = 8'h5D;
		16'h6FA3: out_word = 8'h32;
		16'h6FA4: out_word = 8'h19;
		16'h6FA5: out_word = 8'h5D;
		16'h6FA6: out_word = 8'h32;
		16'h6FA7: out_word = 8'h18;
		16'h6FA8: out_word = 8'h5D;
		16'h6FA9: out_word = 8'h32;
		16'h6FAA: out_word = 8'h0F;
		16'h6FAB: out_word = 8'h5D;
		16'h6FAC: out_word = 8'h32;
		16'h6FAD: out_word = 8'h1F;
		16'h6FAE: out_word = 8'h5D;
		16'h6FAF: out_word = 8'h3E;
		16'h6FB0: out_word = 8'hFF;
		16'h6FB1: out_word = 8'hD3;
		16'h6FB2: out_word = 8'hFF;
		16'h6FB3: out_word = 8'h32;
		16'h6FB4: out_word = 8'h3A;
		16'h6FB5: out_word = 8'h5C;
		16'h6FB6: out_word = 8'h32;
		16'h6FB7: out_word = 8'h16;
		16'h6FB8: out_word = 8'h5D;
		16'h6FB9: out_word = 8'h32;
		16'h6FBA: out_word = 8'h0C;
		16'h6FBB: out_word = 8'h5D;
		16'h6FBC: out_word = 8'h3E;
		16'h6FBD: out_word = 8'hC9;
		16'h6FBE: out_word = 8'h32;
		16'h6FBF: out_word = 8'hC2;
		16'h6FC0: out_word = 8'h5C;
		16'h6FC1: out_word = 8'h3E;
		16'h6FC2: out_word = 8'hD0;
		16'h6FC3: out_word = 8'hD3;
		16'h6FC4: out_word = 8'h1F;
		16'h6FC5: out_word = 8'hC9;
		16'h6FC6: out_word = 8'hCD;
		16'h6FC7: out_word = 8'h0C;
		16'h6FC8: out_word = 8'h05;
		16'h6FC9: out_word = 8'h7E;
		16'h6FCA: out_word = 8'hB7;
		16'h6FCB: out_word = 8'hCA;
		16'h6FCC: out_word = 8'hAC;
		16'h6FCD: out_word = 8'h03;
		16'h6FCE: out_word = 8'hFE;
		16'h6FCF: out_word = 8'h01;
		16'h6FD0: out_word = 8'hCC;
		16'h6FD1: out_word = 8'h07;
		16'h6FD2: out_word = 8'h05;
		16'h6FD3: out_word = 8'hC0;
		16'h6FD4: out_word = 8'h18;
		16'h6FD5: out_word = 8'hF0;
		16'h6FD6: out_word = 8'h06;
		16'h6FD7: out_word = 8'h01;
		16'h6FD8: out_word = 8'h21;
		16'h6FD9: out_word = 8'h25;
		16'h6FDA: out_word = 8'h5D;
		16'h6FDB: out_word = 8'hC3;
		16'h6FDC: out_word = 8'h67;
		16'h6FDD: out_word = 8'h1E;
		16'h6FDE: out_word = 8'hE5;
		16'h6FDF: out_word = 8'hED;
		16'h6FE0: out_word = 8'h5B;
		16'h6FE1: out_word = 8'hF4;
		16'h6FE2: out_word = 8'h5C;
		16'h6FE3: out_word = 8'hCD;
		16'h6FE4: out_word = 8'hD6;
		16'h6FE5: out_word = 8'h2F;
		16'h6FE6: out_word = 8'h3A;
		16'h6FE7: out_word = 8'hDB;
		16'h6FE8: out_word = 8'h5C;
		16'h6FE9: out_word = 8'hD1;
		16'h6FEA: out_word = 8'hB7;
		16'h6FEB: out_word = 8'hC8;
		16'h6FEC: out_word = 8'h4F;
		16'h6FED: out_word = 8'h21;
		16'h6FEE: out_word = 8'h25;
		16'h6FEF: out_word = 8'h5D;
		16'h6FF0: out_word = 8'hED;
		16'h6FF1: out_word = 8'hB0;
		16'h6FF2: out_word = 8'hC9;
		16'h6FF3: out_word = 8'hCF;
		16'h6FF4: out_word = 8'h2A;
		16'h6FF5: out_word = 8'hD0;
		16'h6FF6: out_word = 8'hD1;
		16'h6FF7: out_word = 8'hE6;
		16'h6FF8: out_word = 8'hD2;
		16'h6FF9: out_word = 8'hEF;
		16'h6FFA: out_word = 8'hF8;
		16'h6FFB: out_word = 8'hFE;
		16'h6FFC: out_word = 8'hBE;
		16'h6FFD: out_word = 8'hF4;
		16'h6FFE: out_word = 8'hD5;
		16'h6FFF: out_word = 8'hF7;
		16'h7000: out_word = 8'hD3;
		16'h7001: out_word = 8'hD4;
		16'h7002: out_word = 8'hFF;
		16'h7003: out_word = 8'h34;
		16'h7004: out_word = 8'hEC;
		16'h7005: out_word = 8'h38;
		16'h7006: out_word = 8'hF0;
		16'h7007: out_word = 8'hD6;
		16'h7008: out_word = 8'h33;
		16'h7009: out_word = 8'h04;
		16'h700A: out_word = 8'h18;
		16'h700B: out_word = 8'h10;
		16'h700C: out_word = 8'hC2;
		16'h700D: out_word = 8'h1E;
		16'h700E: out_word = 8'hAB;
		16'h700F: out_word = 8'h16;
		16'h7010: out_word = 8'h3A;
		16'h7011: out_word = 8'h05;
		16'h7012: out_word = 8'h87;
		16'h7013: out_word = 8'h07;
		16'h7014: out_word = 8'h15;
		16'h7015: out_word = 8'h18;
		16'h7016: out_word = 8'hD0;
		16'h7017: out_word = 8'h1A;
		16'h7018: out_word = 8'hFB;
		16'h7019: out_word = 8'h1C;
		16'h701A: out_word = 8'hA5;
		16'h701B: out_word = 8'h19;
		16'h701C: out_word = 8'hA9;
		16'h701D: out_word = 8'h19;
		16'h701E: out_word = 8'hB1;
		16'h701F: out_word = 8'h19;
		16'h7020: out_word = 8'h4D;
		16'h7021: out_word = 8'h1D;
		16'h7022: out_word = 8'h82;
		16'h7023: out_word = 8'h21;
		16'h7024: out_word = 8'h56;
		16'h7025: out_word = 8'h26;
		16'h7026: out_word = 8'h90;
		16'h7027: out_word = 8'h06;
		16'h7028: out_word = 8'hFD;
		16'h7029: out_word = 8'h31;
		16'h702A: out_word = 8'hA1;
		16'h702B: out_word = 8'h2D;
		16'h702C: out_word = 8'hDB;
		16'h702D: out_word = 8'h3A;
		16'h702E: out_word = 8'hCE;
		16'h702F: out_word = 8'h11;
		16'h7030: out_word = 8'h10;
		16'h7031: out_word = 8'h18;
		16'h7032: out_word = 8'h2A;
		16'h7033: out_word = 8'h59;
		16'h7034: out_word = 8'h5C;
		16'h7035: out_word = 8'h22;
		16'h7036: out_word = 8'h11;
		16'h7037: out_word = 8'h5D;
		16'h7038: out_word = 8'h22;
		16'h7039: out_word = 8'hD9;
		16'h703A: out_word = 8'h5C;
		16'h703B: out_word = 8'h3E;
		16'h703C: out_word = 8'hFF;
		16'h703D: out_word = 8'h32;
		16'h703E: out_word = 8'hD6;
		16'h703F: out_word = 8'h5C;
		16'h7040: out_word = 8'h21;
		16'h7041: out_word = 8'hDB;
		16'h7042: out_word = 8'h5C;
		16'h7043: out_word = 8'h22;
		16'h7044: out_word = 8'hD7;
		16'h7045: out_word = 8'h5C;
		16'h7046: out_word = 8'h18;
		16'h7047: out_word = 8'h0F;
		16'h7048: out_word = 8'h22;
		16'h7049: out_word = 8'h11;
		16'h704A: out_word = 8'h5D;
		16'h704B: out_word = 8'h22;
		16'h704C: out_word = 8'hD9;
		16'h704D: out_word = 8'h5C;
		16'h704E: out_word = 8'hCD;
		16'h704F: out_word = 8'hE1;
		16'h7050: out_word = 8'h30;
		16'h7051: out_word = 8'hC0;
		16'h7052: out_word = 8'h23;
		16'h7053: out_word = 8'h23;
		16'h7054: out_word = 8'h22;
		16'h7055: out_word = 8'hD7;
		16'h7056: out_word = 8'h5C;
		16'h7057: out_word = 8'hCD;
		16'h7058: out_word = 8'hA9;
		16'h7059: out_word = 8'h30;
		16'h705A: out_word = 8'h20;
		16'h705B: out_word = 8'h2B;
		16'h705C: out_word = 8'hEB;
		16'h705D: out_word = 8'h13;
		16'h705E: out_word = 8'h06;
		16'h705F: out_word = 8'h00;
		16'h7060: out_word = 8'h21;
		16'h7061: out_word = 8'hC8;
		16'h7062: out_word = 8'h31;
		16'h7063: out_word = 8'h09;
		16'h7064: out_word = 8'h7E;
		16'h7065: out_word = 8'h2A;
		16'h7066: out_word = 8'hD9;
		16'h7067: out_word = 8'h5C;
		16'h7068: out_word = 8'h77;
		16'h7069: out_word = 8'h23;
		16'h706A: out_word = 8'hEB;
		16'h706B: out_word = 8'hE7;
		16'h706C: out_word = 8'hDD;
		16'h706D: out_word = 8'h19;
		16'h706E: out_word = 8'hC5;
		16'h706F: out_word = 8'hE7;
		16'h7070: out_word = 8'hE8;
		16'h7071: out_word = 8'h19;
		16'h7072: out_word = 8'hC1;
		16'h7073: out_word = 8'h3A;
		16'h7074: out_word = 8'hD6;
		16'h7075: out_word = 8'h5C;
		16'h7076: out_word = 8'hB7;
		16'h7077: out_word = 8'h20;
		16'h7078: out_word = 8'h0E;
		16'h7079: out_word = 8'h2A;
		16'h707A: out_word = 8'hD7;
		16'h707B: out_word = 8'h5C;
		16'h707C: out_word = 8'h5E;
		16'h707D: out_word = 8'h23;
		16'h707E: out_word = 8'h56;
		16'h707F: out_word = 8'hEB;
		16'h7080: out_word = 8'hB7;
		16'h7081: out_word = 8'hED;
		16'h7082: out_word = 8'h42;
		16'h7083: out_word = 8'hEB;
		16'h7084: out_word = 8'h72;
		16'h7085: out_word = 8'h2B;
		16'h7086: out_word = 8'h73;
		16'h7087: out_word = 8'h2A;
		16'h7088: out_word = 8'hD9;
		16'h7089: out_word = 8'h5C;
		16'h708A: out_word = 8'h7E;
		16'h708B: out_word = 8'hFE;
		16'h708C: out_word = 8'h0D;
		16'h708D: out_word = 8'hC8;
		16'h708E: out_word = 8'h23;
		16'h708F: out_word = 8'h22;
		16'h7090: out_word = 8'hD9;
		16'h7091: out_word = 8'h5C;
		16'h7092: out_word = 8'h7E;
		16'h7093: out_word = 8'hFE;
		16'h7094: out_word = 8'h0D;
		16'h7095: out_word = 8'hC8;
		16'h7096: out_word = 8'hFE;
		16'h7097: out_word = 8'h22;
		16'h7098: out_word = 8'h20;
		16'h7099: out_word = 8'hBD;
		16'h709A: out_word = 8'h23;
		16'h709B: out_word = 8'h7E;
		16'h709C: out_word = 8'hFE;
		16'h709D: out_word = 8'h0D;
		16'h709E: out_word = 8'hC8;
		16'h709F: out_word = 8'hFE;
		16'h70A0: out_word = 8'h22;
		16'h70A1: out_word = 8'h20;
		16'h70A2: out_word = 8'hF7;
		16'h70A3: out_word = 8'h23;
		16'h70A4: out_word = 8'h22;
		16'h70A5: out_word = 8'hD9;
		16'h70A6: out_word = 8'h5C;
		16'h70A7: out_word = 8'h18;
		16'h70A8: out_word = 8'hAE;
		16'h70A9: out_word = 8'h2A;
		16'h70AA: out_word = 8'hD9;
		16'h70AB: out_word = 8'h5C;
		16'h70AC: out_word = 8'h11;
		16'h70AD: out_word = 8'hFD;
		16'h70AE: out_word = 8'h30;
		16'h70AF: out_word = 8'h0E;
		16'h70B0: out_word = 8'h00;
		16'h70B1: out_word = 8'h7E;
		16'h70B2: out_word = 8'hE6;
		16'h70B3: out_word = 8'hDF;
		16'h70B4: out_word = 8'h47;
		16'h70B5: out_word = 8'hB7;
		16'h70B6: out_word = 8'h20;
		16'h70B7: out_word = 8'h03;
		16'h70B8: out_word = 8'h23;
		16'h70B9: out_word = 8'h18;
		16'h70BA: out_word = 8'hF6;
		16'h70BB: out_word = 8'h1A;
		16'h70BC: out_word = 8'hE6;
		16'h70BD: out_word = 8'h80;
		16'h70BE: out_word = 8'h20;
		16'h70BF: out_word = 8'h08;
		16'h70C0: out_word = 8'h1A;
		16'h70C1: out_word = 8'hB8;
		16'h70C2: out_word = 8'h20;
		16'h70C3: out_word = 8'h15;
		16'h70C4: out_word = 8'h23;
		16'h70C5: out_word = 8'h13;
		16'h70C6: out_word = 8'h18;
		16'h70C7: out_word = 8'hE9;
		16'h70C8: out_word = 8'h1A;
		16'h70C9: out_word = 8'hE6;
		16'h70CA: out_word = 8'h7F;
		16'h70CB: out_word = 8'hB8;
		16'h70CC: out_word = 8'hC8;
		16'h70CD: out_word = 8'h0C;
		16'h70CE: out_word = 8'h2A;
		16'h70CF: out_word = 8'hD9;
		16'h70D0: out_word = 8'h5C;
		16'h70D1: out_word = 8'h13;
		16'h70D2: out_word = 8'h1A;
		16'h70D3: out_word = 8'hFE;
		16'h70D4: out_word = 8'hFF;
		16'h70D5: out_word = 8'h20;
		16'h70D6: out_word = 8'hDA;
		16'h70D7: out_word = 8'hB7;
		16'h70D8: out_word = 8'hC9;
		16'h70D9: out_word = 8'h13;
		16'h70DA: out_word = 8'h1A;
		16'h70DB: out_word = 8'hE6;
		16'h70DC: out_word = 8'h80;
		16'h70DD: out_word = 8'h28;
		16'h70DE: out_word = 8'hFA;
		16'h70DF: out_word = 8'h18;
		16'h70E0: out_word = 8'hEC;
		16'h70E1: out_word = 8'h2A;
		16'h70E2: out_word = 8'h45;
		16'h70E3: out_word = 8'h5C;
		16'h70E4: out_word = 8'h23;
		16'h70E5: out_word = 8'h23;
		16'h70E6: out_word = 8'h7C;
		16'h70E7: out_word = 8'hB5;
		16'h70E8: out_word = 8'h28;
		16'h70E9: out_word = 8'h0A;
		16'h70EA: out_word = 8'hAF;
		16'h70EB: out_word = 8'h32;
		16'h70EC: out_word = 8'hD6;
		16'h70ED: out_word = 8'h5C;
		16'h70EE: out_word = 8'h2B;
		16'h70EF: out_word = 8'h2B;
		16'h70F0: out_word = 8'hE7;
		16'h70F1: out_word = 8'h6E;
		16'h70F2: out_word = 8'h19;
		16'h70F3: out_word = 8'hC9;
		16'h70F4: out_word = 8'h3E;
		16'h70F5: out_word = 8'hFF;
		16'h70F6: out_word = 8'h32;
		16'h70F7: out_word = 8'hD6;
		16'h70F8: out_word = 8'h5C;
		16'h70F9: out_word = 8'h2A;
		16'h70FA: out_word = 8'h59;
		16'h70FB: out_word = 8'h5C;
		16'h70FC: out_word = 8'hC9;
		16'h70FD: out_word = 8'h53;
		16'h70FE: out_word = 8'h41;
		16'h70FF: out_word = 8'h56;
		16'h7100: out_word = 8'h45;
		16'h7101: out_word = 8'h80;
		16'h7102: out_word = 8'h53;
		16'h7103: out_word = 8'h41;
		16'h7104: out_word = 8'h56;
		16'h7105: out_word = 8'hC5;
		16'h7106: out_word = 8'h4C;
		16'h7107: out_word = 8'h4F;
		16'h7108: out_word = 8'h41;
		16'h7109: out_word = 8'h44;
		16'h710A: out_word = 8'h80;
		16'h710B: out_word = 8'h4C;
		16'h710C: out_word = 8'h4F;
		16'h710D: out_word = 8'h41;
		16'h710E: out_word = 8'hC4;
		16'h710F: out_word = 8'h52;
		16'h7110: out_word = 8'h55;
		16'h7111: out_word = 8'h4E;
		16'h7112: out_word = 8'h80;
		16'h7113: out_word = 8'h52;
		16'h7114: out_word = 8'h55;
		16'h7115: out_word = 8'hCE;
		16'h7116: out_word = 8'h43;
		16'h7117: out_word = 8'h41;
		16'h7118: out_word = 8'h54;
		16'h7119: out_word = 8'h80;
		16'h711A: out_word = 8'h43;
		16'h711B: out_word = 8'h41;
		16'h711C: out_word = 8'hD4;
		16'h711D: out_word = 8'h45;
		16'h711E: out_word = 8'h52;
		16'h711F: out_word = 8'h41;
		16'h7120: out_word = 8'h53;
		16'h7121: out_word = 8'h45;
		16'h7122: out_word = 8'h80;
		16'h7123: out_word = 8'h45;
		16'h7124: out_word = 8'h52;
		16'h7125: out_word = 8'h41;
		16'h7126: out_word = 8'h53;
		16'h7127: out_word = 8'hC5;
		16'h7128: out_word = 8'h4E;
		16'h7129: out_word = 8'h45;
		16'h712A: out_word = 8'h57;
		16'h712B: out_word = 8'h80;
		16'h712C: out_word = 8'h4E;
		16'h712D: out_word = 8'h45;
		16'h712E: out_word = 8'hD7;
		16'h712F: out_word = 8'h4D;
		16'h7130: out_word = 8'h4F;
		16'h7131: out_word = 8'h56;
		16'h7132: out_word = 8'h45;
		16'h7133: out_word = 8'h80;
		16'h7134: out_word = 8'h4D;
		16'h7135: out_word = 8'h4F;
		16'h7136: out_word = 8'h56;
		16'h7137: out_word = 8'hC5;
		16'h7138: out_word = 8'h4D;
		16'h7139: out_word = 8'h45;
		16'h713A: out_word = 8'h52;
		16'h713B: out_word = 8'h47;
		16'h713C: out_word = 8'h45;
		16'h713D: out_word = 8'h80;
		16'h713E: out_word = 8'h4D;
		16'h713F: out_word = 8'h45;
		16'h7140: out_word = 8'h52;
		16'h7141: out_word = 8'h47;
		16'h7142: out_word = 8'hC5;
		16'h7143: out_word = 8'h50;
		16'h7144: out_word = 8'h45;
		16'h7145: out_word = 8'h45;
		16'h7146: out_word = 8'h4B;
		16'h7147: out_word = 8'h80;
		16'h7148: out_word = 8'h50;
		16'h7149: out_word = 8'h45;
		16'h714A: out_word = 8'h45;
		16'h714B: out_word = 8'hCB;
		16'h714C: out_word = 8'h50;
		16'h714D: out_word = 8'h4F;
		16'h714E: out_word = 8'h4B;
		16'h714F: out_word = 8'h45;
		16'h7150: out_word = 8'h80;
		16'h7151: out_word = 8'h50;
		16'h7152: out_word = 8'h4F;
		16'h7153: out_word = 8'h4B;
		16'h7154: out_word = 8'hC5;
		16'h7155: out_word = 8'h4F;
		16'h7156: out_word = 8'h50;
		16'h7157: out_word = 8'h45;
		16'h7158: out_word = 8'h4E;
		16'h7159: out_word = 8'h83;
		16'h715A: out_word = 8'h43;
		16'h715B: out_word = 8'h4C;
		16'h715C: out_word = 8'h4F;
		16'h715D: out_word = 8'h53;
		16'h715E: out_word = 8'h45;
		16'h715F: out_word = 8'h83;
		16'h7160: out_word = 8'h43;
		16'h7161: out_word = 8'h4F;
		16'h7162: out_word = 8'h44;
		16'h7163: out_word = 8'h45;
		16'h7164: out_word = 8'h80;
		16'h7165: out_word = 8'h43;
		16'h7166: out_word = 8'h4F;
		16'h7167: out_word = 8'h44;
		16'h7168: out_word = 8'hC5;
		16'h7169: out_word = 8'h52;
		16'h716A: out_word = 8'h4E;
		16'h716B: out_word = 8'h44;
		16'h716C: out_word = 8'h80;
		16'h716D: out_word = 8'h52;
		16'h716E: out_word = 8'h4E;
		16'h716F: out_word = 8'hC4;
		16'h7170: out_word = 8'h44;
		16'h7171: out_word = 8'h41;
		16'h7172: out_word = 8'h54;
		16'h7173: out_word = 8'h41;
		16'h7174: out_word = 8'h80;
		16'h7175: out_word = 8'h44;
		16'h7176: out_word = 8'h41;
		16'h7177: out_word = 8'h54;
		16'h7178: out_word = 8'hC1;
		16'h7179: out_word = 8'h53;
		16'h717A: out_word = 8'h43;
		16'h717B: out_word = 8'h52;
		16'h717C: out_word = 8'h45;
		16'h717D: out_word = 8'h45;
		16'h717E: out_word = 8'h4E;
		16'h717F: out_word = 8'h04;
		16'h7180: out_word = 8'h84;
		16'h7181: out_word = 8'h53;
		16'h7182: out_word = 8'h43;
		16'h7183: out_word = 8'h52;
		16'h7184: out_word = 8'h45;
		16'h7185: out_word = 8'h45;
		16'h7186: out_word = 8'h4E;
		16'h7187: out_word = 8'h84;
		16'h7188: out_word = 8'h43;
		16'h7189: out_word = 8'h4F;
		16'h718A: out_word = 8'h50;
		16'h718B: out_word = 8'h59;
		16'h718C: out_word = 8'h80;
		16'h718D: out_word = 8'h43;
		16'h718E: out_word = 8'h4F;
		16'h718F: out_word = 8'h50;
		16'h7190: out_word = 8'hD9;
		16'h7191: out_word = 8'h46;
		16'h7192: out_word = 8'h4F;
		16'h7193: out_word = 8'h52;
		16'h7194: out_word = 8'h4D;
		16'h7195: out_word = 8'h41;
		16'h7196: out_word = 8'h54;
		16'h7197: out_word = 8'h80;
		16'h7198: out_word = 8'h46;
		16'h7199: out_word = 8'h4F;
		16'h719A: out_word = 8'h52;
		16'h719B: out_word = 8'h4D;
		16'h719C: out_word = 8'h41;
		16'h719D: out_word = 8'hD4;
		16'h719E: out_word = 8'h47;
		16'h719F: out_word = 8'h4F;
		16'h71A0: out_word = 8'h54;
		16'h71A1: out_word = 8'h4F;
		16'h71A2: out_word = 8'h80;
		16'h71A3: out_word = 8'h47;
		16'h71A4: out_word = 8'h4F;
		16'h71A5: out_word = 8'h54;
		16'h71A6: out_word = 8'hCF;
		16'h71A7: out_word = 8'h4C;
		16'h71A8: out_word = 8'h49;
		16'h71A9: out_word = 8'h53;
		16'h71AA: out_word = 8'h54;
		16'h71AB: out_word = 8'h80;
		16'h71AC: out_word = 8'h4C;
		16'h71AD: out_word = 8'h49;
		16'h71AE: out_word = 8'h53;
		16'h71AF: out_word = 8'hD4;
		16'h71B0: out_word = 8'h4C;
		16'h71B1: out_word = 8'h49;
		16'h71B2: out_word = 8'h4E;
		16'h71B3: out_word = 8'h45;
		16'h71B4: out_word = 8'h80;
		16'h71B5: out_word = 8'h4C;
		16'h71B6: out_word = 8'h49;
		16'h71B7: out_word = 8'h4E;
		16'h71B8: out_word = 8'hC5;
		16'h71B9: out_word = 8'h56;
		16'h71BA: out_word = 8'h45;
		16'h71BB: out_word = 8'h52;
		16'h71BC: out_word = 8'h49;
		16'h71BD: out_word = 8'h46;
		16'h71BE: out_word = 8'h59;
		16'h71BF: out_word = 8'h80;
		16'h71C0: out_word = 8'h56;
		16'h71C1: out_word = 8'h45;
		16'h71C2: out_word = 8'h52;
		16'h71C3: out_word = 8'h49;
		16'h71C4: out_word = 8'h46;
		16'h71C5: out_word = 8'hD9;
		16'h71C6: out_word = 8'hFF;
		16'h71C7: out_word = 8'hFF;
		16'h71C8: out_word = 8'hF8;
		16'h71C9: out_word = 8'hF8;
		16'h71CA: out_word = 8'hEF;
		16'h71CB: out_word = 8'hEF;
		16'h71CC: out_word = 8'hF7;
		16'h71CD: out_word = 8'hF7;
		16'h71CE: out_word = 8'hCF;
		16'h71CF: out_word = 8'hCF;
		16'h71D0: out_word = 8'hD2;
		16'h71D1: out_word = 8'hD2;
		16'h71D2: out_word = 8'hE6;
		16'h71D3: out_word = 8'hE6;
		16'h71D4: out_word = 8'hD1;
		16'h71D5: out_word = 8'hD1;
		16'h71D6: out_word = 8'hD5;
		16'h71D7: out_word = 8'hD5;
		16'h71D8: out_word = 8'hBE;
		16'h71D9: out_word = 8'hBE;
		16'h71DA: out_word = 8'hF4;
		16'h71DB: out_word = 8'hF4;
		16'h71DC: out_word = 8'hD3;
		16'h71DD: out_word = 8'hD4;
		16'h71DE: out_word = 8'hAF;
		16'h71DF: out_word = 8'hAF;
		16'h71E0: out_word = 8'hA5;
		16'h71E1: out_word = 8'hA5;
		16'h71E2: out_word = 8'hE4;
		16'h71E3: out_word = 8'hE4;
		16'h71E4: out_word = 8'hAA;
		16'h71E5: out_word = 8'hAA;
		16'h71E6: out_word = 8'hFF;
		16'h71E7: out_word = 8'hFF;
		16'h71E8: out_word = 8'hD0;
		16'h71E9: out_word = 8'hD0;
		16'h71EA: out_word = 8'hEC;
		16'h71EB: out_word = 8'hEC;
		16'h71EC: out_word = 8'hF0;
		16'h71ED: out_word = 8'hF0;
		16'h71EE: out_word = 8'hCA;
		16'h71EF: out_word = 8'hCA;
		16'h71F0: out_word = 8'hD6;
		16'h71F1: out_word = 8'hD6;
		16'h71F2: out_word = 8'h00;
		16'h71F3: out_word = 8'h2A;
		16'h71F4: out_word = 8'h4F;
		16'h71F5: out_word = 8'h5C;
		16'h71F6: out_word = 8'hB7;
		16'h71F7: out_word = 8'h01;
		16'h71F8: out_word = 8'h25;
		16'h71F9: out_word = 8'h5D;
		16'h71FA: out_word = 8'hED;
		16'h71FB: out_word = 8'h42;
		16'h71FC: out_word = 8'hC9;
		16'h71FD: out_word = 8'hCD;
		16'h71FE: out_word = 8'h03;
		16'h71FF: out_word = 8'h32;
		16'h7200: out_word = 8'hC3;
		16'h7201: out_word = 8'hE1;
		16'h7202: out_word = 8'h03;
		16'h7203: out_word = 8'h3E;
		16'h7204: out_word = 8'hD7;
		16'h7205: out_word = 8'h01;
		16'h7206: out_word = 8'hFD;
		16'h7207: out_word = 8'h7F;
		16'h7208: out_word = 8'hED;
		16'h7209: out_word = 8'h79;
		16'h720A: out_word = 8'h32;
		16'h720B: out_word = 8'h00;
		16'h720C: out_word = 8'hC0;
		16'h720D: out_word = 8'h32;
		16'h720E: out_word = 8'hF0;
		16'h720F: out_word = 8'hFF;
		16'h7210: out_word = 8'h3E;
		16'h7211: out_word = 8'h10;
		16'h7212: out_word = 8'hED;
		16'h7213: out_word = 8'h79;
		16'h7214: out_word = 8'hC9;
		16'h7215: out_word = 8'hFF;
		16'h7216: out_word = 8'hFF;
		16'h7217: out_word = 8'hFF;
		16'h7218: out_word = 8'hFF;
		16'h7219: out_word = 8'hFF;
		16'h721A: out_word = 8'hFF;
		16'h721B: out_word = 8'hFF;
		16'h721C: out_word = 8'h3E;
		16'h721D: out_word = 8'h0D;
		16'h721E: out_word = 8'h32;
		16'h721F: out_word = 8'h20;
		16'h7220: out_word = 8'h5D;
		16'h7221: out_word = 8'hC3;
		16'h7222: out_word = 8'h1D;
		16'h7223: out_word = 8'h02;
		16'h7224: out_word = 8'hE5;
		16'h7225: out_word = 8'hC5;
		16'h7226: out_word = 8'hF5;
		16'h7227: out_word = 8'hD5;
		16'h7228: out_word = 8'h3E;
		16'h7229: out_word = 8'hED;
		16'h722A: out_word = 8'h32;
		16'h722B: out_word = 8'h86;
		16'h722C: out_word = 8'h5C;
		16'h722D: out_word = 8'h3E;
		16'h722E: out_word = 8'h0C;
		16'h722F: out_word = 8'h32;
		16'h7230: out_word = 8'h8A;
		16'h7231: out_word = 8'h5C;
		16'h7232: out_word = 8'h7B;
		16'h7233: out_word = 8'h18;
		16'h7234: out_word = 8'h08;
		16'h7235: out_word = 8'h7E;
		16'h7236: out_word = 8'hFE;
		16'h7237: out_word = 8'hFF;
		16'h7238: out_word = 8'hC8;
		16'h7239: out_word = 8'hD7;
		16'h723A: out_word = 8'h23;
		16'h723B: out_word = 8'h18;
		16'h723C: out_word = 8'hF8;
		16'h723D: out_word = 8'h06;
		16'h723E: out_word = 8'h30;
		16'h723F: out_word = 8'hD6;
		16'h7240: out_word = 8'h0A;
		16'h7241: out_word = 8'h38;
		16'h7242: out_word = 8'h03;
		16'h7243: out_word = 8'h04;
		16'h7244: out_word = 8'h18;
		16'h7245: out_word = 8'hF9;
		16'h7246: out_word = 8'hF5;
		16'h7247: out_word = 8'h78;
		16'h7248: out_word = 8'hD7;
		16'h7249: out_word = 8'hF1;
		16'h724A: out_word = 8'hC6;
		16'h724B: out_word = 8'h3A;
		16'h724C: out_word = 8'hD7;
		16'h724D: out_word = 8'hD1;
		16'h724E: out_word = 8'hF1;
		16'h724F: out_word = 8'hC1;
		16'h7250: out_word = 8'hE1;
		16'h7251: out_word = 8'hFB;
		16'h7252: out_word = 8'hC3;
		16'h7253: out_word = 8'h44;
		16'h7254: out_word = 8'h3E;
		16'h7255: out_word = 8'hFF;
		16'h7256: out_word = 8'hFF;
		16'h7257: out_word = 8'hFF;
		16'h7258: out_word = 8'h46;
		16'h7259: out_word = 8'h6F;
		16'h725A: out_word = 8'h72;
		16'h725B: out_word = 8'h6D;
		16'h725C: out_word = 8'h61;
		16'h725D: out_word = 8'h74;
		16'h725E: out_word = 8'h20;
		16'h725F: out_word = 8'h74;
		16'h7260: out_word = 8'h72;
		16'h7261: out_word = 8'h61;
		16'h7262: out_word = 8'h63;
		16'h7263: out_word = 8'h6B;
		16'h7264: out_word = 8'h20;
		16'h7265: out_word = 8'h20;
		16'h7266: out_word = 8'h20;
		16'h7267: out_word = 8'h20;
		16'h7268: out_word = 8'h20;
		16'h7269: out_word = 8'h20;
		16'h726A: out_word = 8'h20;
		16'h726B: out_word = 8'h53;
		16'h726C: out_word = 8'h69;
		16'h726D: out_word = 8'h64;
		16'h726E: out_word = 8'h65;
		16'h726F: out_word = 8'h00;
		16'h7270: out_word = 8'hFF;
		16'h7271: out_word = 8'hFF;
		16'h7272: out_word = 8'hFF;
		16'h7273: out_word = 8'h16;
		16'h7274: out_word = 8'h00;
		16'h7275: out_word = 8'h00;
		16'h7276: out_word = 8'h46;
		16'h7277: out_word = 8'h69;
		16'h7278: out_word = 8'h6C;
		16'h7279: out_word = 8'h65;
		16'h727A: out_word = 8'h20;
		16'h727B: out_word = 8'h22;
		16'h727C: out_word = 8'h13;
		16'h727D: out_word = 8'h01;
		16'h727E: out_word = 8'hFF;
		16'h727F: out_word = 8'h13;
		16'h7280: out_word = 8'h00;
		16'h7281: out_word = 8'h22;
		16'h7282: out_word = 8'h0D;
		16'h7283: out_word = 8'h45;
		16'h7284: out_word = 8'h78;
		16'h7285: out_word = 8'h69;
		16'h7286: out_word = 8'h73;
		16'h7287: out_word = 8'h74;
		16'h7288: out_word = 8'h73;
		16'h7289: out_word = 8'h21;
		16'h728A: out_word = 8'h4F;
		16'h728B: out_word = 8'h76;
		16'h728C: out_word = 8'h65;
		16'h728D: out_word = 8'h72;
		16'h728E: out_word = 8'h77;
		16'h728F: out_word = 8'h72;
		16'h7290: out_word = 8'h69;
		16'h7291: out_word = 8'h74;
		16'h7292: out_word = 8'h65;
		16'h7293: out_word = 8'h3F;
		16'h7294: out_word = 8'h28;
		16'h7295: out_word = 8'h59;
		16'h7296: out_word = 8'h2F;
		16'h7297: out_word = 8'h4E;
		16'h7298: out_word = 8'h2F;
		16'h7299: out_word = 8'h41;
		16'h729A: out_word = 8'h64;
		16'h729B: out_word = 8'h64;
		16'h729C: out_word = 8'h29;
		16'h729D: out_word = 8'hFF;
		16'h729E: out_word = 8'h43;
		16'h729F: out_word = 8'h6F;
		16'h72A0: out_word = 8'h6D;
		16'h72A1: out_word = 8'h70;
		16'h72A2: out_word = 8'h6C;
		16'h72A3: out_word = 8'h65;
		16'h72A4: out_word = 8'h74;
		16'h72A5: out_word = 8'h65;
		16'h72A6: out_word = 8'h0D;
		16'h72A7: out_word = 8'h4E;
		16'h72A8: out_word = 8'h61;
		16'h72A9: out_word = 8'h6D;
		16'h72AA: out_word = 8'h65;
		16'h72AB: out_word = 8'h3A;
		16'h72AC: out_word = 8'h00;
		16'h72AD: out_word = 8'h46;
		16'h72AE: out_word = 8'h4F;
		16'h72AF: out_word = 8'h52;
		16'h72B0: out_word = 8'h4D;
		16'h72B1: out_word = 8'h41;
		16'h72B2: out_word = 8'h54;
		16'h72B3: out_word = 8'h3A;
		16'h72B4: out_word = 8'h20;
		16'h72B5: out_word = 8'h20;
		16'h72B6: out_word = 8'h20;
		16'h72B7: out_word = 8'h31;
		16'h72B8: out_word = 8'h20;
		16'h72B9: out_word = 8'h2D;
		16'h72BA: out_word = 8'h20;
		16'h72BB: out_word = 8'h4E;
		16'h72BC: out_word = 8'h6F;
		16'h72BD: out_word = 8'h72;
		16'h72BE: out_word = 8'h6D;
		16'h72BF: out_word = 8'h61;
		16'h72C0: out_word = 8'h6C;
		16'h72C1: out_word = 8'h20;
		16'h72C2: out_word = 8'h20;
		16'h72C3: out_word = 8'h20;
		16'h72C4: out_word = 8'h0D;
		16'h72C5: out_word = 8'h17;
		16'h72C6: out_word = 8'h0A;
		16'h72C7: out_word = 8'h20;
		16'h72C8: out_word = 8'h32;
		16'h72C9: out_word = 8'h20;
		16'h72CA: out_word = 8'h2D;
		16'h72CB: out_word = 8'h20;
		16'h72CC: out_word = 8'h54;
		16'h72CD: out_word = 8'h75;
		16'h72CE: out_word = 8'h72;
		16'h72CF: out_word = 8'h62;
		16'h72D0: out_word = 8'h6F;
		16'h72D1: out_word = 8'h0D;
		16'h72D2: out_word = 8'h17;
		16'h72D3: out_word = 8'h0A;
		16'h72D4: out_word = 8'h20;
		16'h72D5: out_word = 8'h33;
		16'h72D6: out_word = 8'h20;
		16'h72D7: out_word = 8'h2D;
		16'h72D8: out_word = 8'h20;
		16'h72D9: out_word = 8'h46;
		16'h72DA: out_word = 8'h61;
		16'h72DB: out_word = 8'h73;
		16'h72DC: out_word = 8'h74;
		16'h72DD: out_word = 8'h20;
		16'h72DE: out_word = 8'h74;
		16'h72DF: out_word = 8'h75;
		16'h72E0: out_word = 8'h72;
		16'h72E1: out_word = 8'h62;
		16'h72E2: out_word = 8'h6F;
		16'h72E3: out_word = 8'h00;
		16'h72E4: out_word = 8'hFF;
		16'h72E5: out_word = 8'hFF;
		16'h72E6: out_word = 8'hFF;
		16'h72E7: out_word = 8'hFF;
		16'h72E8: out_word = 8'hFF;
		16'h72E9: out_word = 8'hFF;
		16'h72EA: out_word = 8'h23;
		16'h72EB: out_word = 8'h3A;
		16'h72EC: out_word = 8'hE8;
		16'h72ED: out_word = 8'h5C;
		16'h72EE: out_word = 8'h77;
		16'h72EF: out_word = 8'hAF;
		16'h72F0: out_word = 8'hC9;
		16'h72F1: out_word = 8'hF5;
		16'h72F2: out_word = 8'h3E;
		16'h72F3: out_word = 8'h31;
		16'h72F4: out_word = 8'h18;
		16'h72F5: out_word = 8'h03;
		16'h72F6: out_word = 8'hF5;
		16'h72F7: out_word = 8'h3E;
		16'h72F8: out_word = 8'h30;
		16'h72F9: out_word = 8'hF5;
		16'h72FA: out_word = 8'h3E;
		16'h72FB: out_word = 8'hF8;
		16'h72FC: out_word = 8'h32;
		16'h72FD: out_word = 8'h86;
		16'h72FE: out_word = 8'h5C;
		16'h72FF: out_word = 8'h3E;
		16'h7300: out_word = 8'h17;
		16'h7301: out_word = 8'h32;
		16'h7302: out_word = 8'h8A;
		16'h7303: out_word = 8'h5C;
		16'h7304: out_word = 8'hF1;
		16'h7305: out_word = 8'hD7;
		16'h7306: out_word = 8'hF1;
		16'h7307: out_word = 8'hC3;
		16'h7308: out_word = 8'hFD;
		16'h7309: out_word = 8'h1F;
		16'h730A: out_word = 8'hCD;
		16'h730B: out_word = 8'h9F;
		16'h730C: out_word = 8'h1D;
		16'h730D: out_word = 8'h21;
		16'h730E: out_word = 8'h73;
		16'h730F: out_word = 8'h32;
		16'h7310: out_word = 8'hCD;
		16'h7311: out_word = 8'h35;
		16'h7312: out_word = 8'h32;
		16'h7313: out_word = 8'hCD;
		16'h7314: out_word = 8'h29;
		16'h7315: out_word = 8'h33;
		16'h7316: out_word = 8'h21;
		16'h7317: out_word = 8'h7F;
		16'h7318: out_word = 8'h32;
		16'h7319: out_word = 8'hCD;
		16'h731A: out_word = 8'h35;
		16'h731B: out_word = 8'h32;
		16'h731C: out_word = 8'h21;
		16'h731D: out_word = 8'h00;
		16'h731E: out_word = 8'h40;
		16'h731F: out_word = 8'h2B;
		16'h7320: out_word = 8'h7C;
		16'h7321: out_word = 8'hB5;
		16'h7322: out_word = 8'h20;
		16'h7323: out_word = 8'hFB;
		16'h7324: out_word = 8'hCD;
		16'h7325: out_word = 8'h52;
		16'h7326: out_word = 8'h10;
		16'h7327: out_word = 8'h18;
		16'h7328: out_word = 8'h0F;
		16'h7329: out_word = 8'h3A;
		16'h732A: out_word = 8'hF6;
		16'h732B: out_word = 8'h5C;
		16'h732C: out_word = 8'hC6;
		16'h732D: out_word = 8'h41;
		16'h732E: out_word = 8'hD7;
		16'h732F: out_word = 8'h3E;
		16'h7330: out_word = 8'h3A;
		16'h7331: out_word = 8'hD7;
		16'h7332: out_word = 8'h21;
		16'h7333: out_word = 8'hDD;
		16'h7334: out_word = 8'h5C;
		16'h7335: out_word = 8'hC3;
		16'h7336: out_word = 8'h38;
		16'h7337: out_word = 8'h29;
		16'h7338: out_word = 8'hF5;
		16'h7339: out_word = 8'hCD;
		16'h733A: out_word = 8'h9F;
		16'h733B: out_word = 8'h1D;
		16'h733C: out_word = 8'hF1;
		16'h733D: out_word = 8'hFE;
		16'h733E: out_word = 8'h59;
		16'h733F: out_word = 8'hC8;
		16'h7340: out_word = 8'hFE;
		16'h7341: out_word = 8'h41;
		16'h7342: out_word = 8'hC9;
		16'h7343: out_word = 8'hCD;
		16'h7344: out_word = 8'h5D;
		16'h7345: out_word = 8'h16;
		16'h7346: out_word = 8'h21;
		16'h7347: out_word = 8'hE5;
		16'h7348: out_word = 8'h5C;
		16'h7349: out_word = 8'hCB;
		16'h734A: out_word = 8'hFE;
		16'h734B: out_word = 8'hC9;
		16'h734C: out_word = 8'hCD;
		16'h734D: out_word = 8'h9F;
		16'h734E: out_word = 8'h1D;
		16'h734F: out_word = 8'h21;
		16'h7350: out_word = 8'h58;
		16'h7351: out_word = 8'h32;
		16'h7352: out_word = 8'hDF;
		16'h7353: out_word = 8'hCD;
		16'h7354: out_word = 8'hBD;
		16'h7355: out_word = 8'h20;
		16'h7356: out_word = 8'hCD;
		16'h7357: out_word = 8'h9F;
		16'h7358: out_word = 8'h1D;
		16'h7359: out_word = 8'h21;
		16'h735A: out_word = 8'h9E;
		16'h735B: out_word = 8'h32;
		16'h735C: out_word = 8'hDF;
		16'h735D: out_word = 8'hC9;
		16'h735E: out_word = 8'h50;
		16'h735F: out_word = 8'h72;
		16'h7360: out_word = 8'h65;
		16'h7361: out_word = 8'h73;
		16'h7362: out_word = 8'h73;
		16'h7363: out_word = 8'h20;
		16'h7364: out_word = 8'h52;
		16'h7365: out_word = 8'h20;
		16'h7366: out_word = 8'h74;
		16'h7367: out_word = 8'h6F;
		16'h7368: out_word = 8'h20;
		16'h7369: out_word = 8'h72;
		16'h736A: out_word = 8'h65;
		16'h736B: out_word = 8'h70;
		16'h736C: out_word = 8'h65;
		16'h736D: out_word = 8'h61;
		16'h736E: out_word = 8'h74;
		16'h736F: out_word = 8'hAE;
		16'h7370: out_word = 8'h00;
		16'h7371: out_word = 8'hCD;
		16'h7372: out_word = 8'h9F;
		16'h7373: out_word = 8'h1D;
		16'h7374: out_word = 8'hCD;
		16'h7375: out_word = 8'h11;
		16'h7376: out_word = 8'h3E;
		16'h7377: out_word = 8'hC9;
		16'h7378: out_word = 8'hCD;
		16'h7379: out_word = 8'h9F;
		16'h737A: out_word = 8'h1D;
		16'h737B: out_word = 8'h21;
		16'h737C: out_word = 8'hAD;
		16'h737D: out_word = 8'h32;
		16'h737E: out_word = 8'hDF;
		16'h737F: out_word = 8'hCD;
		16'h7380: out_word = 8'h52;
		16'h7381: out_word = 8'h10;
		16'h7382: out_word = 8'hFE;
		16'h7383: out_word = 8'h11;
		16'h7384: out_word = 8'h28;
		16'h7385: out_word = 8'h0F;
		16'h7386: out_word = 8'hFE;
		16'h7387: out_word = 8'h12;
		16'h7388: out_word = 8'h28;
		16'h7389: out_word = 8'h17;
		16'h738A: out_word = 8'hFE;
		16'h738B: out_word = 8'h13;
		16'h738C: out_word = 8'h28;
		16'h738D: out_word = 8'h18;
		16'h738E: out_word = 8'hFE;
		16'h738F: out_word = 8'h00;
		16'h7390: out_word = 8'hCA;
		16'h7391: out_word = 8'hD3;
		16'h7392: out_word = 8'h01;
		16'h7393: out_word = 8'h18;
		16'h7394: out_word = 8'hEA;
		16'h7395: out_word = 8'h21;
		16'h7396: out_word = 8'hB9;
		16'h7397: out_word = 8'h1F;
		16'h7398: out_word = 8'hAF;
		16'h7399: out_word = 8'h32;
		16'h739A: out_word = 8'hE8;
		16'h739B: out_word = 8'h5C;
		16'h739C: out_word = 8'h22;
		16'h739D: out_word = 8'hE6;
		16'h739E: out_word = 8'h5C;
		16'h739F: out_word = 8'h18;
		16'h73A0: out_word = 8'hD0;
		16'h73A1: out_word = 8'h21;
		16'h73A2: out_word = 8'hAD;
		16'h73A3: out_word = 8'h33;
		16'h73A4: out_word = 8'h18;
		16'h73A5: out_word = 8'hF2;
		16'h73A6: out_word = 8'h3E;
		16'h73A7: out_word = 8'h01;
		16'h73A8: out_word = 8'h21;
		16'h73A9: out_word = 8'hAD;
		16'h73AA: out_word = 8'h33;
		16'h73AB: out_word = 8'h18;
		16'h73AC: out_word = 8'hEC;
		16'h73AD: out_word = 8'h01;
		16'h73AE: out_word = 8'h02;
		16'h73AF: out_word = 8'h03;
		16'h73B0: out_word = 8'h04;
		16'h73B1: out_word = 8'h05;
		16'h73B2: out_word = 8'h06;
		16'h73B3: out_word = 8'h07;
		16'h73B4: out_word = 8'h08;
		16'h73B5: out_word = 8'h09;
		16'h73B6: out_word = 8'h0A;
		16'h73B7: out_word = 8'h0B;
		16'h73B8: out_word = 8'h0C;
		16'h73B9: out_word = 8'h0D;
		16'h73BA: out_word = 8'h0E;
		16'h73BB: out_word = 8'h0F;
		16'h73BC: out_word = 8'h10;
		16'h73BD: out_word = 8'h01;
		16'h73BE: out_word = 8'h7D;
		16'h73BF: out_word = 8'hD6;
		16'h73C0: out_word = 8'h0E;
		16'h73C1: out_word = 8'h6F;
		16'h73C2: out_word = 8'hD0;
		16'h73C3: out_word = 8'h25;
		16'h73C4: out_word = 8'hC9;
		16'h73C5: out_word = 8'hFF;
		16'h73C6: out_word = 8'hFF;
		16'h73C7: out_word = 8'hFF;
		16'h73C8: out_word = 8'hFF;
		16'h73C9: out_word = 8'hFF;
		16'h73CA: out_word = 8'hFF;
		16'h73CB: out_word = 8'hFF;
		16'h73CC: out_word = 8'hFF;
		16'h73CD: out_word = 8'hFF;
		16'h73CE: out_word = 8'h3A;
		16'h73CF: out_word = 8'hE5;
		16'h73D0: out_word = 8'h5C;
		16'h73D1: out_word = 8'hFE;
		16'h73D2: out_word = 8'h42;
		16'h73D3: out_word = 8'h28;
		16'h73D4: out_word = 8'h0D;
		16'h73D5: out_word = 8'hFE;
		16'h73D6: out_word = 8'h44;
		16'h73D7: out_word = 8'h28;
		16'h73D8: out_word = 8'h09;
		16'h73D9: out_word = 8'hFE;
		16'h73DA: out_word = 8'h23;
		16'h73DB: out_word = 8'h28;
		16'h73DC: out_word = 8'h05;
		16'h73DD: out_word = 8'h3E;
		16'h73DE: out_word = 8'h43;
		16'h73DF: out_word = 8'hFF;
		16'h73E0: out_word = 8'hFF;
		16'h73E1: out_word = 8'hFF;
		16'h73E2: out_word = 8'h3A;
		16'h73E3: out_word = 8'hD6;
		16'h73E4: out_word = 8'h5C;
		16'h73E5: out_word = 8'hC9;
		16'h73E6: out_word = 8'hCD;
		16'h73E7: out_word = 8'hF0;
		16'h73E8: out_word = 8'h1C;
		16'h73E9: out_word = 8'hCC;
		16'h73EA: out_word = 8'h43;
		16'h73EB: out_word = 8'h33;
		16'h73EC: out_word = 8'hCD;
		16'h73ED: out_word = 8'h05;
		16'h73EE: out_word = 8'h04;
		16'h73EF: out_word = 8'hCD;
		16'h73F0: out_word = 8'hC4;
		16'h73F1: out_word = 8'h1A;
		16'h73F2: out_word = 8'hC3;
		16'h73F3: out_word = 8'h53;
		16'h73F4: out_word = 8'h1B;
		16'h73F5: out_word = 8'h21;
		16'h73F6: out_word = 8'hE5;
		16'h73F7: out_word = 8'h5C;
		16'h73F8: out_word = 8'hCB;
		16'h73F9: out_word = 8'h7E;
		16'h73FA: out_word = 8'hCB;
		16'h73FB: out_word = 8'hBE;
		16'h73FC: out_word = 8'hCA;
		16'h73FD: out_word = 8'h59;
		16'h73FE: out_word = 8'h1B;
		16'h73FF: out_word = 8'hCD;
		16'h7400: out_word = 8'h0A;
		16'h7401: out_word = 8'h33;
		16'h7402: out_word = 8'hC2;
		16'h7403: out_word = 8'hD3;
		16'h7404: out_word = 8'h01;
		16'h7405: out_word = 8'hFE;
		16'h7406: out_word = 8'h41;
		16'h7407: out_word = 8'hCA;
		16'h7408: out_word = 8'h59;
		16'h7409: out_word = 8'h1B;
		16'h740A: out_word = 8'hED;
		16'h740B: out_word = 8'h5B;
		16'h740C: out_word = 8'hD9;
		16'h740D: out_word = 8'h5C;
		16'h740E: out_word = 8'h1B;
		16'h740F: out_word = 8'h14;
		16'h7410: out_word = 8'h3A;
		16'h7411: out_word = 8'hEA;
		16'h7412: out_word = 8'h5C;
		16'h7413: out_word = 8'hBA;
		16'h7414: out_word = 8'h28;
		16'h7415: out_word = 8'h05;
		16'h7416: out_word = 8'hCD;
		16'h7417: out_word = 8'h26;
		16'h7418: out_word = 8'h29;
		16'h7419: out_word = 8'h18;
		16'h741A: out_word = 8'hD1;
		16'h741B: out_word = 8'h42;
		16'h741C: out_word = 8'h2A;
		16'h741D: out_word = 8'h59;
		16'h741E: out_word = 8'h5C;
		16'h741F: out_word = 8'h36;
		16'h7420: out_word = 8'hAA;
		16'h7421: out_word = 8'h23;
		16'h7422: out_word = 8'hED;
		16'h7423: out_word = 8'h5B;
		16'h7424: out_word = 8'hD1;
		16'h7425: out_word = 8'h5C;
		16'h7426: out_word = 8'h73;
		16'h7427: out_word = 8'h23;
		16'h7428: out_word = 8'h72;
		16'h7429: out_word = 8'h0E;
		16'h742A: out_word = 8'h06;
		16'h742B: out_word = 8'h2A;
		16'h742C: out_word = 8'hDB;
		16'h742D: out_word = 8'h5C;
		16'h742E: out_word = 8'h22;
		16'h742F: out_word = 8'hE8;
		16'h7430: out_word = 8'h5C;
		16'h7431: out_word = 8'h2A;
		16'h7432: out_word = 8'hD7;
		16'h7433: out_word = 8'h5C;
		16'h7434: out_word = 8'h22;
		16'h7435: out_word = 8'hE6;
		16'h7436: out_word = 8'h5C;
		16'h7437: out_word = 8'hED;
		16'h7438: out_word = 8'h5B;
		16'h7439: out_word = 8'hEB;
		16'h743A: out_word = 8'h5C;
		16'h743B: out_word = 8'hCD;
		16'h743C: out_word = 8'h4D;
		16'h743D: out_word = 8'h1E;
		16'h743E: out_word = 8'hED;
		16'h743F: out_word = 8'h4B;
		16'h7440: out_word = 8'h1E;
		16'h7441: out_word = 8'h5D;
		16'h7442: out_word = 8'hCD;
		16'h7443: out_word = 8'hBF;
		16'h7444: out_word = 8'h1B;
		16'h7445: out_word = 8'hCD;
		16'h7446: out_word = 8'h65;
		16'h7447: out_word = 8'h16;
		16'h7448: out_word = 8'hC9;
		16'h7449: out_word = 8'hFB;
		16'h744A: out_word = 8'hC3;
		16'h744B: out_word = 8'h69;
		16'h744C: out_word = 8'h2F;
		16'h744D: out_word = 8'h00;
		16'h744E: out_word = 8'hDD;
		16'h744F: out_word = 8'h7E;
		16'h7450: out_word = 8'h00;
		16'h7451: out_word = 8'hFE;
		16'h7452: out_word = 8'hFF;
		16'h7453: out_word = 8'h20;
		16'h7454: out_word = 8'h06;
		16'h7455: out_word = 8'h3A;
		16'h7456: out_word = 8'h6F;
		16'h7457: out_word = 8'hF8;
		16'h7458: out_word = 8'hDD;
		16'h7459: out_word = 8'h77;
		16'h745A: out_word = 8'h00;
		16'h745B: out_word = 8'hCD;
		16'h745C: out_word = 8'hFA;
		16'h745D: out_word = 8'hF7;
		16'h745E: out_word = 8'hCD;
		16'h745F: out_word = 8'h16;
		16'h7460: out_word = 8'hF8;
		16'h7461: out_word = 8'hC3;
		16'h7462: out_word = 8'h46;
		16'h7463: out_word = 8'hF6;
		16'h7464: out_word = 8'hCD;
		16'h7465: out_word = 8'h70;
		16'h7466: out_word = 8'hF8;
		16'h7467: out_word = 8'hCD;
		16'h7468: out_word = 8'h26;
		16'h7469: out_word = 8'hF8;
		16'h746A: out_word = 8'hDD;
		16'h746B: out_word = 8'h34;
		16'h746C: out_word = 8'h00;
		16'h746D: out_word = 8'h3A;
		16'h746E: out_word = 8'h6F;
		16'h746F: out_word = 8'hF8;
		16'h7470: out_word = 8'h3C;
		16'h7471: out_word = 8'hDD;
		16'h7472: out_word = 8'hBE;
		16'h7473: out_word = 8'h00;
		16'h7474: out_word = 8'hDD;
		16'h7475: out_word = 8'h7E;
		16'h7476: out_word = 8'h00;
		16'h7477: out_word = 8'h20;
		16'h7478: out_word = 8'h04;
		16'h7479: out_word = 8'hAF;
		16'h747A: out_word = 8'hDD;
		16'h747B: out_word = 8'h77;
		16'h747C: out_word = 8'h00;
		16'h747D: out_word = 8'hCD;
		16'h747E: out_word = 8'hFA;
		16'h747F: out_word = 8'hF7;
		16'h7480: out_word = 8'hCD;
		16'h7481: out_word = 8'h16;
		16'h7482: out_word = 8'hF8;
		16'h7483: out_word = 8'hC3;
		16'h7484: out_word = 8'h46;
		16'h7485: out_word = 8'hF6;
		16'h7486: out_word = 8'hCD;
		16'h7487: out_word = 8'h70;
		16'h7488: out_word = 8'hF8;
		16'h7489: out_word = 8'hCD;
		16'h748A: out_word = 8'h26;
		16'h748B: out_word = 8'hF8;
		16'h748C: out_word = 8'hDD;
		16'h748D: out_word = 8'h35;
		16'h748E: out_word = 8'h00;
		16'h748F: out_word = 8'hDD;
		16'h7490: out_word = 8'h35;
		16'h7491: out_word = 8'h00;
		16'h7492: out_word = 8'hDD;
		16'h7493: out_word = 8'h35;
		16'h7494: out_word = 8'h00;
		16'h7495: out_word = 8'hDD;
		16'h7496: out_word = 8'hCB;
		16'h7497: out_word = 8'h00;
		16'h7498: out_word = 8'h7E;
		16'h7499: out_word = 8'hDD;
		16'h749A: out_word = 8'h7E;
		16'h749B: out_word = 8'h00;
		16'h749C: out_word = 8'h28;
		16'h749D: out_word = 8'h15;
		16'h749E: out_word = 8'h06;
		16'h749F: out_word = 8'h03;
		16'h74A0: out_word = 8'h80;
		16'h74A1: out_word = 8'h47;
		16'h74A2: out_word = 8'hC5;
		16'h74A3: out_word = 8'h3A;
		16'h74A4: out_word = 8'h6F;
		16'h74A5: out_word = 8'hF8;
		16'h74A6: out_word = 8'h90;
		16'h74A7: out_word = 8'h38;
		16'h74A8: out_word = 8'h03;
		16'h74A9: out_word = 8'hF1;
		16'h74AA: out_word = 8'h18;
		16'h74AB: out_word = 8'hF2;
		16'h74AC: out_word = 8'hF1;
		16'h74AD: out_word = 8'h3D;
		16'h74AE: out_word = 8'h3D;
		16'h74AF: out_word = 8'h3D;
		16'h74B0: out_word = 8'hDD;
		16'h74B1: out_word = 8'h77;
		16'h74B2: out_word = 8'h00;
		16'h74B3: out_word = 8'hCD;
		16'h74B4: out_word = 8'hFA;
		16'h74B5: out_word = 8'hF7;
		16'h74B6: out_word = 8'hCD;
		16'h74B7: out_word = 8'h16;
		16'h74B8: out_word = 8'hF8;
		16'h74B9: out_word = 8'hC3;
		16'h74BA: out_word = 8'h46;
		16'h74BB: out_word = 8'hF6;
		16'h74BC: out_word = 8'hCD;
		16'h74BD: out_word = 8'h70;
		16'h74BE: out_word = 8'hF8;
		16'h74BF: out_word = 8'hCD;
		16'h74C0: out_word = 8'h26;
		16'h74C1: out_word = 8'hF8;
		16'h74C2: out_word = 8'hDD;
		16'h74C3: out_word = 8'h34;
		16'h74C4: out_word = 8'h00;
		16'h74C5: out_word = 8'hDD;
		16'h74C6: out_word = 8'h34;
		16'h74C7: out_word = 8'h00;
		16'h74C8: out_word = 8'hDD;
		16'h74C9: out_word = 8'h34;
		16'h74CA: out_word = 8'h00;
		16'h74CB: out_word = 8'h3A;
		16'h74CC: out_word = 8'h6F;
		16'h74CD: out_word = 8'hF8;
		16'h74CE: out_word = 8'hDD;
		16'h74CF: out_word = 8'h9E;
		16'h74D0: out_word = 8'h00;
		16'h74D1: out_word = 8'hDD;
		16'h74D2: out_word = 8'h7E;
		16'h74D3: out_word = 8'h00;
		16'h74D4: out_word = 8'h30;
		16'h74D5: out_word = 8'h0B;
		16'h74D6: out_word = 8'h06;
		16'h74D7: out_word = 8'h03;
		16'h74D8: out_word = 8'h90;
		16'h74D9: out_word = 8'h30;
		16'h74DA: out_word = 8'hFD;
		16'h74DB: out_word = 8'h3C;
		16'h74DC: out_word = 8'h3C;
		16'h74DD: out_word = 8'h3C;
		16'h74DE: out_word = 8'hDD;
		16'h74DF: out_word = 8'h77;
		16'h74E0: out_word = 8'h00;
		16'h74E1: out_word = 8'hCD;
		16'h74E2: out_word = 8'hFA;
		16'h74E3: out_word = 8'hF7;
		16'h74E4: out_word = 8'hCD;
		16'h74E5: out_word = 8'h16;
		16'h74E6: out_word = 8'hF8;
		16'h74E7: out_word = 8'hC3;
		16'h74E8: out_word = 8'h46;
		16'h74E9: out_word = 8'hF6;
		16'h74EA: out_word = 8'hCD;
		16'h74EB: out_word = 8'h6B;
		16'h74EC: out_word = 8'h0D;
		16'h74ED: out_word = 8'h3E;
		16'h74EE: out_word = 8'h03;
		16'h74EF: out_word = 8'hCD;
		16'h74F0: out_word = 8'hCB;
		16'h74F1: out_word = 8'hF8;
		16'h74F2: out_word = 8'hC3;
		16'h74F3: out_word = 8'h56;
		16'h74F4: out_word = 8'hF5;
		16'h74F5: out_word = 8'h01;
		16'h74F6: out_word = 8'hFD;
		16'h74F7: out_word = 8'hFF;
		16'h74F8: out_word = 8'h3E;
		16'h74F9: out_word = 8'h07;
		16'h74FA: out_word = 8'hED;
		16'h74FB: out_word = 8'h79;
		16'h74FC: out_word = 8'h06;
		16'h74FD: out_word = 8'hBF;
		16'h74FE: out_word = 8'h3E;
		16'h74FF: out_word = 8'hFF;
		16'h7500: out_word = 8'hED;
		16'h7501: out_word = 8'h79;
		16'h7502: out_word = 8'hCD;
		16'h7503: out_word = 8'h70;
		16'h7504: out_word = 8'hF8;
		16'h7505: out_word = 8'h3E;
		16'h7506: out_word = 8'h07;
		16'h7507: out_word = 8'h32;
		16'h7508: out_word = 8'h48;
		16'h7509: out_word = 8'h5C;
		16'h750A: out_word = 8'h32;
		16'h750B: out_word = 8'h8D;
		16'h750C: out_word = 8'h5C;
		16'h750D: out_word = 8'h2F;
		16'h750E: out_word = 8'h32;
		16'h750F: out_word = 8'h3B;
		16'h7510: out_word = 8'h5D;
		16'h7511: out_word = 8'h21;
		16'h7512: out_word = 8'h00;
		16'h7513: out_word = 8'h3C;
		16'h7514: out_word = 8'h22;
		16'h7515: out_word = 8'h36;
		16'h7516: out_word = 8'h5C;
		16'h7517: out_word = 8'hDD;
		16'h7518: out_word = 8'h6E;
		16'h7519: out_word = 8'h00;
		16'h751A: out_word = 8'h26;
		16'h751B: out_word = 8'h00;
		16'h751C: out_word = 8'h29;
		16'h751D: out_word = 8'h29;
		16'h751E: out_word = 8'h29;
		16'h751F: out_word = 8'h11;
		16'h7520: out_word = 8'h00;
		16'h7521: out_word = 8'hA0;
		16'h7522: out_word = 8'h19;
		16'h7523: out_word = 8'h11;
		16'h7524: out_word = 8'hF0;
		16'h7525: out_word = 8'hF7;
		16'h7526: out_word = 8'h01;
		16'h7527: out_word = 8'h08;
		16'h7528: out_word = 8'h00;
		16'h7529: out_word = 8'hED;
		16'h752A: out_word = 8'hB0;
		16'h752B: out_word = 8'h2A;
		16'h752C: out_word = 8'h32;
		16'h752D: out_word = 8'hF6;
		16'h752E: out_word = 8'h22;
		16'h752F: out_word = 8'h3D;
		16'h7530: out_word = 8'h5C;
		16'h7531: out_word = 8'h21;
		16'h7532: out_word = 8'hEC;
		16'h7533: out_word = 8'hF7;
		16'h7534: out_word = 8'h22;
		16'h7535: out_word = 8'h5D;
		16'h7536: out_word = 8'h5C;
		16'h7537: out_word = 8'hCD;
		16'h7538: out_word = 8'h6B;
		16'h7539: out_word = 8'h0D;
		16'h753A: out_word = 8'hF3;
		16'h753B: out_word = 8'hE1;
		16'h753C: out_word = 8'hD9;
		16'h753D: out_word = 8'hC1;
		16'h753E: out_word = 8'hD1;
		16'h753F: out_word = 8'hE1;
		16'h7540: out_word = 8'hF1;
		16'h7541: out_word = 8'hCD;
		16'h7542: out_word = 8'h03;
		16'h7543: out_word = 8'h3D;
		16'h7544: out_word = 8'hEA;
		16'h7545: out_word = 8'h3A;
		16'h7546: out_word = 8'hF7;
		16'h7547: out_word = 8'h22;
		16'h7548: out_word = 8'h62;
		16'h7549: out_word = 8'h6F;
		16'h754A: out_word = 8'h6F;
		16'h754B: out_word = 8'h74;
		16'h754C: out_word = 8'h20;
		16'h754D: out_word = 8'h20;
		16'h754E: out_word = 8'h20;
		16'h754F: out_word = 8'h20;
		16'h7550: out_word = 8'h22;
		16'h7551: out_word = 8'h0D;
		16'h7552: out_word = 8'hD5;
		16'h7553: out_word = 8'h3C;
		16'h7554: out_word = 8'h21;
		16'h7555: out_word = 8'h02;
		16'h7556: out_word = 8'h58;
		16'h7557: out_word = 8'h11;
		16'h7558: out_word = 8'h0A;
		16'h7559: out_word = 8'h00;
		16'h755A: out_word = 8'h3D;
		16'h755B: out_word = 8'h28;
		16'h755C: out_word = 8'h0F;
		16'h755D: out_word = 8'h19;
		16'h755E: out_word = 8'h3D;
		16'h755F: out_word = 8'h28;
		16'h7560: out_word = 8'h0B;
		16'h7561: out_word = 8'h19;
		16'h7562: out_word = 8'h3D;
		16'h7563: out_word = 8'h28;
		16'h7564: out_word = 8'h07;
		16'h7565: out_word = 8'h13;
		16'h7566: out_word = 8'h13;
		16'h7567: out_word = 8'h19;
		16'h7568: out_word = 8'h1B;
		16'h7569: out_word = 8'h1B;
		16'h756A: out_word = 8'h18;
		16'h756B: out_word = 8'hEE;
		16'h756C: out_word = 8'hD1;
		16'h756D: out_word = 8'hC9;
		16'h756E: out_word = 8'hE5;
		16'h756F: out_word = 8'hD9;
		16'h7570: out_word = 8'hE1;
		16'h7571: out_word = 8'h3E;
		16'h7572: out_word = 8'h70;
		16'h7573: out_word = 8'hE5;
		16'h7574: out_word = 8'hD1;
		16'h7575: out_word = 8'h13;
		16'h7576: out_word = 8'h01;
		16'h7577: out_word = 8'h07;
		16'h7578: out_word = 8'h00;
		16'h7579: out_word = 8'h77;
		16'h757A: out_word = 8'hED;
		16'h757B: out_word = 8'hB0;
		16'h757C: out_word = 8'hD9;
		16'h757D: out_word = 8'hC9;
		16'h757E: out_word = 8'hE5;
		16'h757F: out_word = 8'hD9;
		16'h7580: out_word = 8'hE1;
		16'h7581: out_word = 8'h3E;
		16'h7582: out_word = 8'h42;
		16'h7583: out_word = 8'hE5;
		16'h7584: out_word = 8'hD1;
		16'h7585: out_word = 8'h13;
		16'h7586: out_word = 8'h01;
		16'h7587: out_word = 8'h07;
		16'h7588: out_word = 8'h00;
		16'h7589: out_word = 8'h77;
		16'h758A: out_word = 8'hED;
		16'h758B: out_word = 8'hB0;
		16'h758C: out_word = 8'hD9;
		16'h758D: out_word = 8'hC9;
		16'h758E: out_word = 8'hE5;
		16'h758F: out_word = 8'hD5;
		16'h7590: out_word = 8'hED;
		16'h7591: out_word = 8'h52;
		16'h7592: out_word = 8'h7E;
		16'h7593: out_word = 8'h06;
		16'h7594: out_word = 8'h20;
		16'h7595: out_word = 8'h98;
		16'h7596: out_word = 8'h38;
		16'h7597: out_word = 8'h2B;
		16'h7598: out_word = 8'hDD;
		16'h7599: out_word = 8'h21;
		16'h759A: out_word = 8'h81;
		16'h759B: out_word = 8'hF9;
		16'h759C: out_word = 8'hE5;
		16'h759D: out_word = 8'h01;
		16'h759E: out_word = 8'h00;
		16'h759F: out_word = 8'h08;
		16'h75A0: out_word = 8'h7E;
		16'h75A1: out_word = 8'hDD;
		16'h75A2: out_word = 8'hBE;
		16'h75A3: out_word = 8'h00;
		16'h75A4: out_word = 8'h20;
		16'h75A5: out_word = 8'h01;
		16'h75A6: out_word = 8'h0C;
		16'h75A7: out_word = 8'h23;
		16'h75A8: out_word = 8'hDD;
		16'h75A9: out_word = 8'h23;
		16'h75AA: out_word = 8'h10;
		16'h75AB: out_word = 8'hF4;
		16'h75AC: out_word = 8'h79;
		16'h75AD: out_word = 8'hFE;
		16'h75AE: out_word = 8'h08;
		16'h75AF: out_word = 8'h20;
		16'h75B0: out_word = 8'h03;
		16'h75B1: out_word = 8'hE1;
		16'h75B2: out_word = 8'h18;
		16'h75B3: out_word = 8'h0F;
		16'h75B4: out_word = 8'hD9;
		16'h75B5: out_word = 8'hE1;
		16'h75B6: out_word = 8'h01;
		16'h75B7: out_word = 8'h08;
		16'h75B8: out_word = 8'h00;
		16'h75B9: out_word = 8'hED;
		16'h75BA: out_word = 8'hB0;
		16'h75BB: out_word = 8'hD9;
		16'h75BC: out_word = 8'h3A;
		16'h75BD: out_word = 8'h6E;
		16'h75BE: out_word = 8'hF8;
		16'h75BF: out_word = 8'h3C;
		16'h75C0: out_word = 8'h32;
		16'h75C1: out_word = 8'h6E;
		16'h75C2: out_word = 8'hF8;
		16'h75C3: out_word = 8'hD1;
		16'h75C4: out_word = 8'hE1;
		16'h75C5: out_word = 8'hC9;
		16'h75C6: out_word = 8'h00;
		16'h75C7: out_word = 8'h00;
		16'h75C8: out_word = 8'hF5;
		16'h75C9: out_word = 8'hC5;
		16'h75CA: out_word = 8'h06;
		16'h75CB: out_word = 8'hD2;
		16'h75CC: out_word = 8'hC5;
		16'h75CD: out_word = 8'hAF;
		16'h75CE: out_word = 8'hD3;
		16'h75CF: out_word = 8'hFE;
		16'h75D0: out_word = 8'hCB;
		16'h75D1: out_word = 8'h18;
		16'h75D2: out_word = 8'h10;
		16'h75D3: out_word = 8'hFE;
		16'h75D4: out_word = 8'hCB;
		16'h75D5: out_word = 8'hE7;
		16'h75D6: out_word = 8'hD3;
		16'h75D7: out_word = 8'hFE;
		16'h75D8: out_word = 8'hC1;
		16'h75D9: out_word = 8'h05;
		16'h75DA: out_word = 8'h10;
		16'h75DB: out_word = 8'hF0;
		16'h75DC: out_word = 8'hC1;
		16'h75DD: out_word = 8'hF1;
		16'h75DE: out_word = 8'hC9;
		16'h75DF: out_word = 8'hAF;
		16'h75E0: out_word = 8'hFD;
		16'h75E1: out_word = 8'hBE;
		16'h75E2: out_word = 8'h47;
		16'h75E3: out_word = 8'hC2;
		16'h75E4: out_word = 8'h56;
		16'h75E5: out_word = 8'hF5;
		16'h75E6: out_word = 8'hCD;
		16'h75E7: out_word = 8'h6E;
		16'h75E8: out_word = 8'h0D;
		16'h75E9: out_word = 8'h3E;
		16'h75EA: out_word = 8'h02;
		16'h75EB: out_word = 8'hCD;
		16'h75EC: out_word = 8'h01;
		16'h75ED: out_word = 8'h16;
		16'h75EE: out_word = 8'hAF;
		16'h75EF: out_word = 8'hCD;
		16'h75F0: out_word = 8'hCB;
		16'h75F1: out_word = 8'hF8;
		16'h75F2: out_word = 8'h3E;
		16'h75F3: out_word = 8'h01;
		16'h75F4: out_word = 8'hCD;
		16'h75F5: out_word = 8'h01;
		16'h75F6: out_word = 8'h16;
		16'h75F7: out_word = 8'hFD;
		16'h75F8: out_word = 8'h36;
		16'h75F9: out_word = 8'h47;
		16'h75FA: out_word = 8'hFE;
		16'h75FB: out_word = 8'hC3;
		16'h75FC: out_word = 8'h95;
		16'h75FD: out_word = 8'hF7;
		16'h75FE: out_word = 8'hAF;
		16'h75FF: out_word = 8'hFD;
		16'h7600: out_word = 8'hBE;
		16'h7601: out_word = 8'h47;
		16'h7602: out_word = 8'hC2;
		16'h7603: out_word = 8'h56;
		16'h7604: out_word = 8'hF5;
		16'h7605: out_word = 8'hCD;
		16'h7606: out_word = 8'h6E;
		16'h7607: out_word = 8'h0D;
		16'h7608: out_word = 8'h3E;
		16'h7609: out_word = 8'h02;
		16'h760A: out_word = 8'hCD;
		16'h760B: out_word = 8'h01;
		16'h760C: out_word = 8'h16;
		16'h760D: out_word = 8'h3E;
		16'h760E: out_word = 8'h01;
		16'h760F: out_word = 8'hCD;
		16'h7610: out_word = 8'hCB;
		16'h7611: out_word = 8'hF8;
		16'h7612: out_word = 8'h3E;
		16'h7613: out_word = 8'h3F;
		16'h7614: out_word = 8'h32;
		16'h7615: out_word = 8'h6E;
		16'h7616: out_word = 8'hF8;
		16'h7617: out_word = 8'h01;
		16'h7618: out_word = 8'hFF;
		16'h7619: out_word = 8'hFF;
		16'h761A: out_word = 8'h00;
		16'h761B: out_word = 8'h10;
		16'h761C: out_word = 8'hFD;
		16'h761D: out_word = 8'h0D;
		16'h761E: out_word = 8'h20;
		16'h761F: out_word = 8'hFA;
		16'h7620: out_word = 8'hC3;
		16'h7621: out_word = 8'hB4;
		16'h7622: out_word = 8'hF5;
		16'h7623: out_word = 8'h11;
		16'h7624: out_word = 8'hD1;
		16'h7625: out_word = 8'hF8;
		16'h7626: out_word = 8'hC3;
		16'h7627: out_word = 8'h0A;
		16'h7628: out_word = 8'h0C;
		16'h7629: out_word = 8'h80;
		16'h762A: out_word = 8'h16;
		16'h762B: out_word = 8'h0A;
		16'h762C: out_word = 8'h05;
		16'h762D: out_word = 8'h21;
		16'h762E: out_word = 8'h21;
		16'h762F: out_word = 8'h21;
		16'h7630: out_word = 8'h20;
		16'h7631: out_word = 8'h4E;
		16'h7632: out_word = 8'h4F;
		16'h7633: out_word = 8'h20;
		16'h7634: out_word = 8'h20;
		16'h7635: out_word = 8'h50;
		16'h7636: out_word = 8'h52;
		16'h7637: out_word = 8'h4F;
		16'h7638: out_word = 8'h47;
		16'h7639: out_word = 8'h52;
		16'h763A: out_word = 8'h41;
		16'h763B: out_word = 8'h4D;
		16'h763C: out_word = 8'h53;
		16'h763D: out_word = 8'h20;
		16'h763E: out_word = 8'h21;
		16'h763F: out_word = 8'h21;
		16'h7640: out_word = 8'h21;
		16'h7641: out_word = 8'hA0;
		16'h7642: out_word = 8'h16;
		16'h7643: out_word = 8'h0A;
		16'h7644: out_word = 8'h03;
		16'h7645: out_word = 8'h10;
		16'h7646: out_word = 8'h04;
		16'h7647: out_word = 8'h4D;
		16'h7648: out_word = 8'h4F;
		16'h7649: out_word = 8'h52;
		16'h764A: out_word = 8'h45;
		16'h764B: out_word = 8'h20;
		16'h764C: out_word = 8'h54;
		16'h764D: out_word = 8'h48;
		16'h764E: out_word = 8'h41;
		16'h764F: out_word = 8'h4E;
		16'h7650: out_word = 8'h20;
		16'h7651: out_word = 8'h36;
		16'h7652: out_word = 8'h33;
		16'h7653: out_word = 8'h20;
		16'h7654: out_word = 8'h42;
		16'h7655: out_word = 8'h41;
		16'h7656: out_word = 8'h53;
		16'h7657: out_word = 8'h49;
		16'h7658: out_word = 8'h43;
		16'h7659: out_word = 8'h20;
		16'h765A: out_word = 8'h46;
		16'h765B: out_word = 8'h49;
		16'h765C: out_word = 8'h4C;
		16'h765D: out_word = 8'h45;
		16'h765E: out_word = 8'h53;
		16'h765F: out_word = 8'hA0;
		16'h7660: out_word = 8'h11;
		16'h7661: out_word = 8'h00;
		16'h7662: out_word = 8'h10;
		16'h7663: out_word = 8'h04;
		16'h7664: out_word = 8'h13;
		16'h7665: out_word = 8'h01;
		16'h7666: out_word = 8'h20;
		16'h7667: out_word = 8'h20;
		16'h7668: out_word = 8'h20;
		16'h7669: out_word = 8'h20;
		16'h766A: out_word = 8'h20;
		16'h766B: out_word = 8'h2D;
		16'h766C: out_word = 8'h3D;
		16'h766D: out_word = 8'h4E;
		16'h766E: out_word = 8'h65;
		16'h766F: out_word = 8'h77;
		16'h7670: out_word = 8'h20;
		16'h7671: out_word = 8'h52;
		16'h7672: out_word = 8'h4F;
		16'h7673: out_word = 8'h4D;
		16'h7674: out_word = 8'h20;
		16'h7675: out_word = 8'h62;
		16'h7676: out_word = 8'h6F;
		16'h7677: out_word = 8'h6F;
		16'h7678: out_word = 8'h74;
		16'h7679: out_word = 8'h20;
		16'h767A: out_word = 8'h76;
		16'h767B: out_word = 8'h31;
		16'h767C: out_word = 8'h2E;
		16'h767D: out_word = 8'h30;
		16'h767E: out_word = 8'h36;
		16'h767F: out_word = 8'h3D;
		16'h7680: out_word = 8'h2D;
		16'h7681: out_word = 8'h06;
		16'h7682: out_word = 8'h52;
		16'h7683: out_word = 8'h65;
		16'h7684: out_word = 8'h6D;
		16'h7685: out_word = 8'h69;
		16'h7686: out_word = 8'h78;
		16'h7687: out_word = 8'h20;
		16'h7688: out_word = 8'h62;
		16'h7689: out_word = 8'h79;
		16'h768A: out_word = 8'h20;
		16'h768B: out_word = 8'h43;
		16'h768C: out_word = 8'h6F;
		16'h768D: out_word = 8'h6D;
		16'h768E: out_word = 8'h70;
		16'h768F: out_word = 8'h6F;
		16'h7690: out_word = 8'h57;
		16'h7691: out_word = 8'h65;
		16'h7692: out_word = 8'h6C;
		16'h7693: out_word = 8'h6C;
		16'h7694: out_word = 8'h63;
		16'h7695: out_word = 8'h6F;
		16'h7696: out_word = 8'h6D;
		16'h7697: out_word = 8'h65;
		16'h7698: out_word = 8'h20;
		16'h7699: out_word = 8'h30;
		16'h769A: out_word = 8'h35;
		16'h769B: out_word = 8'h2E;
		16'h769C: out_word = 8'h30;
		16'h769D: out_word = 8'h32;
		16'h769E: out_word = 8'h2E;
		16'h769F: out_word = 8'h39;
		16'h76A0: out_word = 8'h39;
		16'h76A1: out_word = 8'hAE;
		16'h76A2: out_word = 8'h10;
		16'h76A3: out_word = 8'h02;
		16'h76A4: out_word = 8'h13;
		16'h76A5: out_word = 8'h01;
		16'h76A6: out_word = 8'h20;
		16'h76A7: out_word = 8'h20;
		16'h76A8: out_word = 8'h20;
		16'h76A9: out_word = 8'h20;
		16'h76AA: out_word = 8'h20;
		16'h76AB: out_word = 8'h20;
		16'h76AC: out_word = 8'h20;
		16'h76AD: out_word = 8'h49;
		16'h76AE: out_word = 8'h4E;
		16'h76AF: out_word = 8'h53;
		16'h76B0: out_word = 8'h45;
		16'h76B1: out_word = 8'h52;
		16'h76B2: out_word = 8'h54;
		16'h76B3: out_word = 8'h20;
		16'h76B4: out_word = 8'h4E;
		16'h76B5: out_word = 8'h45;
		16'h76B6: out_word = 8'h57;
		16'h76B7: out_word = 8'h20;
		16'h76B8: out_word = 8'h44;
		16'h76B9: out_word = 8'h49;
		16'h76BA: out_word = 8'h53;
		16'h76BB: out_word = 8'h4B;
		16'h76BC: out_word = 8'h06;
		16'h76BD: out_word = 8'h20;
		16'h76BE: out_word = 8'h20;
		16'h76BF: out_word = 8'h20;
		16'h76C0: out_word = 8'h20;
		16'h76C1: out_word = 8'h20;
		16'h76C2: out_word = 8'h46;
		16'h76C3: out_word = 8'h4F;
		16'h76C4: out_word = 8'h52;
		16'h76C5: out_word = 8'h20;
		16'h76C6: out_word = 8'h52;
		16'h76C7: out_word = 8'h45;
		16'h76C8: out_word = 8'h41;
		16'h76C9: out_word = 8'h44;
		16'h76CA: out_word = 8'h49;
		16'h76CB: out_word = 8'h4E;
		16'h76CC: out_word = 8'h47;
		16'h76CD: out_word = 8'h20;
		16'h76CE: out_word = 8'h43;
		16'h76CF: out_word = 8'h41;
		16'h76D0: out_word = 8'h54;
		16'h76D1: out_word = 8'h41;
		16'h76D2: out_word = 8'h4C;
		16'h76D3: out_word = 8'h4F;
		16'h76D4: out_word = 8'h47;
		16'h76D5: out_word = 8'h55;
		16'h76D6: out_word = 8'h45;
		16'h76D7: out_word = 8'h2E;
		16'h76D8: out_word = 8'hA0;
		16'h76D9: out_word = 8'h62;
		16'h76DA: out_word = 8'h6F;
		16'h76DB: out_word = 8'h6F;
		16'h76DC: out_word = 8'h74;
		16'h76DD: out_word = 8'h20;
		16'h76DE: out_word = 8'h20;
		16'h76DF: out_word = 8'h20;
		16'h76E0: out_word = 8'h20;
		16'h76E1: out_word = 8'h21;
		16'h76E2: out_word = 8'hE1;
		16'h76E3: out_word = 8'h5A;
		16'h76E4: out_word = 8'hE5;
		16'h76E5: out_word = 8'hD1;
		16'h76E6: out_word = 8'h1B;
		16'h76E7: out_word = 8'h01;
		16'h76E8: out_word = 8'h1F;
		16'h76E9: out_word = 8'h00;
		16'h76EA: out_word = 8'hED;
		16'h76EB: out_word = 8'hB0;
		16'h76EC: out_word = 8'h21;
		16'h76ED: out_word = 8'hFF;
		16'h76EE: out_word = 8'h5A;
		16'h76EF: out_word = 8'h3A;
		16'h76F0: out_word = 8'hBA;
		16'h76F1: out_word = 8'hF9;
		16'h76F2: out_word = 8'hB7;
		16'h76F3: out_word = 8'h28;
		16'h76F4: out_word = 8'h0E;
		16'h76F5: out_word = 8'h7E;
		16'h76F6: out_word = 8'hE6;
		16'h76F7: out_word = 8'h07;
		16'h76F8: out_word = 8'h3C;
		16'h76F9: out_word = 8'hFE;
		16'h76FA: out_word = 8'h08;
		16'h76FB: out_word = 8'h20;
		16'h76FC: out_word = 8'h13;
		16'h76FD: out_word = 8'hAF;
		16'h76FE: out_word = 8'h32;
		16'h76FF: out_word = 8'hBA;
		16'h7700: out_word = 8'hF9;
		16'h7701: out_word = 8'h3E;
		16'h7702: out_word = 8'h07;
		16'h7703: out_word = 8'h7E;
		16'h7704: out_word = 8'hE6;
		16'h7705: out_word = 8'h07;
		16'h7706: out_word = 8'h3D;
		16'h7707: out_word = 8'hB7;
		16'h7708: out_word = 8'h20;
		16'h7709: out_word = 8'h06;
		16'h770A: out_word = 8'h2F;
		16'h770B: out_word = 8'h32;
		16'h770C: out_word = 8'hBA;
		16'h770D: out_word = 8'hF9;
		16'h770E: out_word = 8'h3E;
		16'h770F: out_word = 8'h01;
		16'h7710: out_word = 8'h77;
		16'h7711: out_word = 8'hC9;
		16'h7712: out_word = 8'h00;
		16'h7713: out_word = 8'h3E;
		16'h7714: out_word = 8'hC3;
		16'h7715: out_word = 8'h32;
		16'h7716: out_word = 8'hC2;
		16'h7717: out_word = 8'h5C;
		16'h7718: out_word = 8'h21;
		16'h7719: out_word = 8'hE6;
		16'h771A: out_word = 8'hF9;
		16'h771B: out_word = 8'h22;
		16'h771C: out_word = 8'hC3;
		16'h771D: out_word = 8'h5C;
		16'h771E: out_word = 8'hDD;
		16'h771F: out_word = 8'h21;
		16'h7720: out_word = 8'hC1;
		16'h7721: out_word = 8'h2F;
		16'h7722: out_word = 8'hCD;
		16'h7723: out_word = 8'h20;
		16'h7724: out_word = 8'hFA;
		16'h7725: out_word = 8'h3E;
		16'h7726: out_word = 8'h08;
		16'h7727: out_word = 8'h0E;
		16'h7728: out_word = 8'h1F;
		16'h7729: out_word = 8'hDD;
		16'h772A: out_word = 8'h21;
		16'h772B: out_word = 8'h53;
		16'h772C: out_word = 8'h2A;
		16'h772D: out_word = 8'hCD;
		16'h772E: out_word = 8'h20;
		16'h772F: out_word = 8'hFA;
		16'h7730: out_word = 8'hED;
		16'h7731: out_word = 8'h73;
		16'h7732: out_word = 8'hE7;
		16'h7733: out_word = 8'hF9;
		16'h7734: out_word = 8'h11;
		16'h7735: out_word = 8'h00;
		16'h7736: out_word = 8'h00;
		16'h7737: out_word = 8'hDD;
		16'h7738: out_word = 8'h21;
		16'h7739: out_word = 8'h40;
		16'h773A: out_word = 8'h27;
		16'h773B: out_word = 8'hCD;
		16'h773C: out_word = 8'h20;
		16'h773D: out_word = 8'hFA;
		16'h773E: out_word = 8'h31;
		16'h773F: out_word = 8'h00;
		16'h7740: out_word = 8'h00;
		16'h7741: out_word = 8'hDD;
		16'h7742: out_word = 8'h21;
		16'h7743: out_word = 8'hF3;
		16'h7744: out_word = 8'h1F;
		16'h7745: out_word = 8'hCD;
		16'h7746: out_word = 8'h20;
		16'h7747: out_word = 8'hFA;
		16'h7748: out_word = 8'hDD;
		16'h7749: out_word = 8'h21;
		16'h774A: out_word = 8'hEB;
		16'h774B: out_word = 8'h1F;
		16'h774C: out_word = 8'hCD;
		16'h774D: out_word = 8'h20;
		16'h774E: out_word = 8'hFA;
		16'h774F: out_word = 8'hDD;
		16'h7750: out_word = 8'h21;
		16'h7751: out_word = 8'hC1;
		16'h7752: out_word = 8'h2F;
		16'h7753: out_word = 8'hCD;
		16'h7754: out_word = 8'h20;
		16'h7755: out_word = 8'hFA;
		16'h7756: out_word = 8'h3E;
		16'h7757: out_word = 8'hC9;
		16'h7758: out_word = 8'h32;
		16'h7759: out_word = 8'hC2;
		16'h775A: out_word = 8'h5C;
		16'h775B: out_word = 8'h3A;
		16'h775C: out_word = 8'hCD;
		16'h775D: out_word = 8'h5C;
		16'h775E: out_word = 8'hE6;
		16'h775F: out_word = 8'h40;
		16'h7760: out_word = 8'hC9;
		16'h7761: out_word = 8'h3E;
		16'h7762: out_word = 8'h30;
		16'h7763: out_word = 8'h3C;
		16'h7764: out_word = 8'hFE;
		16'h7765: out_word = 8'h33;
		16'h7766: out_word = 8'h32;
		16'h7767: out_word = 8'h0A;
		16'h7768: out_word = 8'hFA;
		16'h7769: out_word = 8'hC2;
		16'h776A: out_word = 8'hD0;
		16'h776B: out_word = 8'hF6;
		16'h776C: out_word = 8'h3E;
		16'h776D: out_word = 8'h30;
		16'h776E: out_word = 8'h32;
		16'h776F: out_word = 8'h0A;
		16'h7770: out_word = 8'hFA;
		16'h7771: out_word = 8'h18;
		16'h7772: out_word = 8'hEE;
		16'h7773: out_word = 8'hF3;
		16'h7774: out_word = 8'hDD;
		16'h7775: out_word = 8'h21;
		16'h7776: out_word = 8'h00;
		16'h7777: out_word = 8'h00;
		16'h7778: out_word = 8'hDD;
		16'h7779: out_word = 8'hE5;
		16'h777A: out_word = 8'hC3;
		16'h777B: out_word = 8'h2F;
		16'h777C: out_word = 8'h3D;
		16'h777D: out_word = 8'hFF;
		16'h777E: out_word = 8'hFF;
		16'h777F: out_word = 8'hFF;
		16'h7780: out_word = 8'hF5;
		16'h7781: out_word = 8'h3A;
		16'h7782: out_word = 8'hCE;
		16'h7783: out_word = 8'h5C;
		16'h7784: out_word = 8'hB7;
		16'h7785: out_word = 8'h28;
		16'h7786: out_word = 8'h0A;
		16'h7787: out_word = 8'hF1;
		16'h7788: out_word = 8'hC5;
		16'h7789: out_word = 8'h47;
		16'h778A: out_word = 8'hDB;
		16'h778B: out_word = 8'h3F;
		16'h778C: out_word = 8'hB8;
		16'h778D: out_word = 8'hC1;
		16'h778E: out_word = 8'hC3;
		16'h778F: out_word = 8'h54;
		16'h7790: out_word = 8'h3E;
		16'h7791: out_word = 8'hF1;
		16'h7792: out_word = 8'hDB;
		16'h7793: out_word = 8'h1F;
		16'h7794: out_word = 8'hE6;
		16'h7795: out_word = 8'h80;
		16'h7796: out_word = 8'hC3;
		16'h7797: out_word = 8'h54;
		16'h7798: out_word = 8'h3E;
		16'h7799: out_word = 8'hFF;
		16'h779A: out_word = 8'h21;
		16'h779B: out_word = 8'hF0;
		16'h779C: out_word = 8'hFF;
		16'h779D: out_word = 8'hAF;
		16'h779E: out_word = 8'hAE;
		16'h779F: out_word = 8'h8C;
		16'h77A0: out_word = 8'h2C;
		16'h77A1: out_word = 8'h20;
		16'h77A2: out_word = 8'hFB;
		16'h77A3: out_word = 8'hFE;
		16'h77A4: out_word = 8'h06;
		16'h77A5: out_word = 8'hCA;
		16'h77A6: out_word = 8'h00;
		16'h77A7: out_word = 8'hC0;
		16'h77A8: out_word = 8'hAF;
		16'h77A9: out_word = 8'hCD;
		16'h77AA: out_word = 8'hC5;
		16'h77AB: out_word = 8'h3C;
		16'h77AC: out_word = 8'h06;
		16'h77AD: out_word = 8'h13;
		16'h77AE: out_word = 8'h26;
		16'h77AF: out_word = 8'h5B;
		16'h77B0: out_word = 8'hAF;
		16'h77B1: out_word = 8'hAE;
		16'h77B2: out_word = 8'h8D;
		16'h77B3: out_word = 8'h8E;
		16'h77B4: out_word = 8'h2C;
		16'h77B5: out_word = 8'h10;
		16'h77B6: out_word = 8'hFA;
		16'h77B7: out_word = 8'hFE;
		16'h77B8: out_word = 8'h68;
		16'h77B9: out_word = 8'hC2;
		16'h77BA: out_word = 8'h4B;
		16'h77BB: out_word = 8'h3C;
		16'h77BC: out_word = 8'hAF;
		16'h77BD: out_word = 8'h32;
		16'h77BE: out_word = 8'h04;
		16'h77BF: out_word = 8'h5B;
		16'h77C0: out_word = 8'h32;
		16'h77C1: out_word = 8'h0D;
		16'h77C2: out_word = 8'h5B;
		16'h77C3: out_word = 8'h21;
		16'h77C4: out_word = 8'hC7;
		16'h77C5: out_word = 8'h00;
		16'h77C6: out_word = 8'h22;
		16'h77C7: out_word = 8'h11;
		16'h77C8: out_word = 8'h5B;
		16'h77C9: out_word = 8'hC3;
		16'h77CA: out_word = 8'h00;
		16'h77CB: out_word = 8'h5B;
		16'h77CC: out_word = 8'hFF;
		16'h77CD: out_word = 8'hE5;
		16'h77CE: out_word = 8'hF5;
		16'h77CF: out_word = 8'hCD;
		16'h77D0: out_word = 8'h08;
		16'h77D1: out_word = 8'h3E;
		16'h77D2: out_word = 8'h47;
		16'h77D3: out_word = 8'hF1;
		16'h77D4: out_word = 8'hE1;
		16'h77D5: out_word = 8'hC3;
		16'h77D6: out_word = 8'h44;
		16'h77D7: out_word = 8'h3E;
		16'h77D8: out_word = 8'h2A;
		16'h77D9: out_word = 8'h11;
		16'h77DA: out_word = 8'h5D;
		16'h77DB: out_word = 8'h23;
		16'h77DC: out_word = 8'h7E;
		16'h77DD: out_word = 8'hFE;
		16'h77DE: out_word = 8'h0D;
		16'h77DF: out_word = 8'h28;
		16'h77E0: out_word = 8'h06;
		16'h77E1: out_word = 8'hCD;
		16'h77E2: out_word = 8'hCD;
		16'h77E3: out_word = 8'h1D;
		16'h77E4: out_word = 8'hC3;
		16'h77E5: out_word = 8'h3D;
		16'h77E6: out_word = 8'h05;
		16'h77E7: out_word = 8'h21;
		16'h77E8: out_word = 8'hEE;
		16'h77E9: out_word = 8'h37;
		16'h77EA: out_word = 8'hDF;
		16'h77EB: out_word = 8'hC3;
		16'h77EC: out_word = 8'hD3;
		16'h77ED: out_word = 8'h01;
		16'h77EE: out_word = 8'h52;
		16'h77EF: out_word = 8'h65;
		16'h77F0: out_word = 8'h6C;
		16'h77F1: out_word = 8'h3A;
		16'h77F2: out_word = 8'h20;
		16'h77F3: out_word = 8'h32;
		16'h77F4: out_word = 8'h32;
		16'h77F5: out_word = 8'h2E;
		16'h77F6: out_word = 8'h30;
		16'h77F7: out_word = 8'h36;
		16'h77F8: out_word = 8'h2E;
		16'h77F9: out_word = 8'h30;
		16'h77FA: out_word = 8'h35;
		16'h77FB: out_word = 8'h0D;
		16'h77FC: out_word = 8'h00;
		16'h77FD: out_word = 8'hFF;
		16'h77FE: out_word = 8'hFF;
		16'h77FF: out_word = 8'hFF;
		16'h7800: out_word = 8'h3A;
		16'h7801: out_word = 8'hF6;
		16'h7802: out_word = 8'h5C;
		16'h7803: out_word = 8'hFE;
		16'h7804: out_word = 8'h03;
		16'h7805: out_word = 8'h28;
		16'h7806: out_word = 8'h09;
		16'h7807: out_word = 8'h3A;
		16'h7808: out_word = 8'hCE;
		16'h7809: out_word = 8'h5C;
		16'h780A: out_word = 8'hCD;
		16'h780B: out_word = 8'h36;
		16'h780C: out_word = 8'h1E;
		16'h780D: out_word = 8'hC3;
		16'h780E: out_word = 8'h70;
		16'h780F: out_word = 8'h1E;
		16'h7810: out_word = 8'hD5;
		16'h7811: out_word = 8'hCD;
		16'h7812: out_word = 8'h37;
		16'h7813: out_word = 8'h38;
		16'h7814: out_word = 8'hC2;
		16'h7815: out_word = 8'hE1;
		16'h7816: out_word = 8'h3E;
		16'h7817: out_word = 8'hD1;
		16'h7818: out_word = 8'hE1;
		16'h7819: out_word = 8'hC1;
		16'h781A: out_word = 8'hAF;
		16'h781B: out_word = 8'hB0;
		16'h781C: out_word = 8'hC8;
		16'h781D: out_word = 8'hC5;
		16'h781E: out_word = 8'hE5;
		16'h781F: out_word = 8'hCD;
		16'h7820: out_word = 8'h80;
		16'h7821: out_word = 8'h38;
		16'h7822: out_word = 8'hE1;
		16'h7823: out_word = 8'h24;
		16'h7824: out_word = 8'hE5;
		16'h7825: out_word = 8'h21;
		16'h7826: out_word = 8'hF4;
		16'h7827: out_word = 8'h5C;
		16'h7828: out_word = 8'h3E;
		16'h7829: out_word = 8'h10;
		16'h782A: out_word = 8'h34;
		16'h782B: out_word = 8'hBE;
		16'h782C: out_word = 8'h20;
		16'h782D: out_word = 8'h04;
		16'h782E: out_word = 8'h36;
		16'h782F: out_word = 8'h00;
		16'h7830: out_word = 8'h23;
		16'h7831: out_word = 8'h34;
		16'h7832: out_word = 8'hE1;
		16'h7833: out_word = 8'hC1;
		16'h7834: out_word = 8'h10;
		16'h7835: out_word = 8'hE7;
		16'h7836: out_word = 8'hC9;
		16'h7837: out_word = 8'hF3;
		16'h7838: out_word = 8'h21;
		16'h7839: out_word = 8'h10;
		16'h783A: out_word = 8'hFF;
		16'h783B: out_word = 8'hCD;
		16'h783C: out_word = 8'h61;
		16'h783D: out_word = 8'h39;
		16'h783E: out_word = 8'hED;
		16'h783F: out_word = 8'h69;
		16'h7840: out_word = 8'h56;
		16'h7841: out_word = 8'h74;
		16'h7842: out_word = 8'h3E;
		16'h7843: out_word = 8'h90;
		16'h7844: out_word = 8'hED;
		16'h7845: out_word = 8'h79;
		16'h7846: out_word = 8'h5E;
		16'h7847: out_word = 8'h75;
		16'h7848: out_word = 8'hED;
		16'h7849: out_word = 8'h69;
		16'h784A: out_word = 8'h44;
		16'h784B: out_word = 8'h78;
		16'h784C: out_word = 8'hBE;
		16'h784D: out_word = 8'h20;
		16'h784E: out_word = 8'h0E;
		16'h784F: out_word = 8'h06;
		16'h7850: out_word = 8'h7F;
		16'h7851: out_word = 8'h72;
		16'h7852: out_word = 8'h3E;
		16'h7853: out_word = 8'h90;
		16'h7854: out_word = 8'hED;
		16'h7855: out_word = 8'h79;
		16'h7856: out_word = 8'h73;
		16'h7857: out_word = 8'hED;
		16'h7858: out_word = 8'h69;
		16'h7859: out_word = 8'h3E;
		16'h785A: out_word = 8'h08;
		16'h785B: out_word = 8'h06;
		16'h785C: out_word = 8'h83;
		16'h785D: out_word = 8'hF5;
		16'h785E: out_word = 8'h32;
		16'h785F: out_word = 8'hFD;
		16'h7860: out_word = 8'h5C;
		16'h7861: out_word = 8'h78;
		16'h7862: out_word = 8'h32;
		16'h7863: out_word = 8'hCB;
		16'h7864: out_word = 8'h5C;
		16'h7865: out_word = 8'hAF;
		16'h7866: out_word = 8'hD3;
		16'h7867: out_word = 8'hFF;
		16'h7868: out_word = 8'h3A;
		16'h7869: out_word = 8'hF6;
		16'h786A: out_word = 8'h5C;
		16'h786B: out_word = 8'hC6;
		16'h786C: out_word = 8'h3C;
		16'h786D: out_word = 8'h32;
		16'h786E: out_word = 8'h16;
		16'h786F: out_word = 8'h5D;
		16'h7870: out_word = 8'hD3;
		16'h7871: out_word = 8'hFF;
		16'h7872: out_word = 8'h3E;
		16'h7873: out_word = 8'hD0;
		16'h7874: out_word = 8'hD3;
		16'h7875: out_word = 8'h1F;
		16'h7876: out_word = 8'h3A;
		16'h7877: out_word = 8'h5C;
		16'h7878: out_word = 8'h5B;
		16'h7879: out_word = 8'h01;
		16'h787A: out_word = 8'hFD;
		16'h787B: out_word = 8'h7F;
		16'h787C: out_word = 8'hED;
		16'h787D: out_word = 8'h79;
		16'h787E: out_word = 8'hF1;
		16'h787F: out_word = 8'hC9;
		16'h7880: out_word = 8'hED;
		16'h7881: out_word = 8'h5B;
		16'h7882: out_word = 8'hF4;
		16'h7883: out_word = 8'h5C;
		16'h7884: out_word = 8'h7C;
		16'h7885: out_word = 8'hFE;
		16'h7886: out_word = 8'hBF;
		16'h7887: out_word = 8'h38;
		16'h7888: out_word = 8'h4B;
		16'h7889: out_word = 8'h3E;
		16'h788A: out_word = 8'hFF;
		16'h788B: out_word = 8'hCD;
		16'h788C: out_word = 8'hA8;
		16'h788D: out_word = 8'h38;
		16'h788E: out_word = 8'h3A;
		16'h788F: out_word = 8'hCE;
		16'h7890: out_word = 8'h5C;
		16'h7891: out_word = 8'hA7;
		16'h7892: out_word = 8'h28;
		16'h7893: out_word = 8'h2E;
		16'h7894: out_word = 8'h11;
		16'h7895: out_word = 8'h25;
		16'h7896: out_word = 8'h5D;
		16'h7897: out_word = 8'h01;
		16'h7898: out_word = 8'h00;
		16'h7899: out_word = 8'h01;
		16'h789A: out_word = 8'hED;
		16'h789B: out_word = 8'hB0;
		16'h789C: out_word = 8'h21;
		16'h789D: out_word = 8'h25;
		16'h789E: out_word = 8'h5D;
		16'h789F: out_word = 8'hED;
		16'h78A0: out_word = 8'h5B;
		16'h78A1: out_word = 8'hF4;
		16'h78A2: out_word = 8'h5C;
		16'h78A3: out_word = 8'hCD;
		16'h78A4: out_word = 8'hD4;
		16'h78A5: out_word = 8'h38;
		16'h78A6: out_word = 8'h3E;
		16'h78A7: out_word = 8'h00;
		16'h78A8: out_word = 8'h08;
		16'h78A9: out_word = 8'h3A;
		16'h78AA: out_word = 8'hCE;
		16'h78AB: out_word = 8'h5C;
		16'h78AC: out_word = 8'h08;
		16'h78AD: out_word = 8'h32;
		16'h78AE: out_word = 8'hCE;
		16'h78AF: out_word = 8'h5C;
		16'h78B0: out_word = 8'hE5;
		16'h78B1: out_word = 8'hD5;
		16'h78B2: out_word = 8'h21;
		16'h78B3: out_word = 8'h25;
		16'h78B4: out_word = 8'h5D;
		16'h78B5: out_word = 8'h11;
		16'h78B6: out_word = 8'h0F;
		16'h78B7: out_word = 8'h00;
		16'h78B8: out_word = 8'hCD;
		16'h78B9: out_word = 8'hD4;
		16'h78BA: out_word = 8'h38;
		16'h78BB: out_word = 8'hD1;
		16'h78BC: out_word = 8'hE1;
		16'h78BD: out_word = 8'h08;
		16'h78BE: out_word = 8'h32;
		16'h78BF: out_word = 8'hCE;
		16'h78C0: out_word = 8'h5C;
		16'h78C1: out_word = 8'hC9;
		16'h78C2: out_word = 8'hE5;
		16'h78C3: out_word = 8'h21;
		16'h78C4: out_word = 8'h25;
		16'h78C5: out_word = 8'h5D;
		16'h78C6: out_word = 8'hCD;
		16'h78C7: out_word = 8'hD4;
		16'h78C8: out_word = 8'h38;
		16'h78C9: out_word = 8'h21;
		16'h78CA: out_word = 8'h25;
		16'h78CB: out_word = 8'h5D;
		16'h78CC: out_word = 8'hD1;
		16'h78CD: out_word = 8'h01;
		16'h78CE: out_word = 8'h00;
		16'h78CF: out_word = 8'h01;
		16'h78D0: out_word = 8'hED;
		16'h78D1: out_word = 8'hB0;
		16'h78D2: out_word = 8'h18;
		16'h78D3: out_word = 8'hD2;
		16'h78D4: out_word = 8'hF3;
		16'h78D5: out_word = 8'hCD;
		16'h78D6: out_word = 8'h61;
		16'h78D7: out_word = 8'h39;
		16'h78D8: out_word = 8'h7A;
		16'h78D9: out_word = 8'h2F;
		16'h78DA: out_word = 8'h0F;
		16'h78DB: out_word = 8'h0F;
		16'h78DC: out_word = 8'hE6;
		16'h78DD: out_word = 8'h3F;
		16'h78DE: out_word = 8'hF5;
		16'h78DF: out_word = 8'hE6;
		16'h78E0: out_word = 8'h27;
		16'h78E1: out_word = 8'hF6;
		16'h78E2: out_word = 8'h10;
		16'h78E3: out_word = 8'h4F;
		16'h78E4: out_word = 8'hF1;
		16'h78E5: out_word = 8'h07;
		16'h78E6: out_word = 8'h07;
		16'h78E7: out_word = 8'h07;
		16'h78E8: out_word = 8'hE6;
		16'h78E9: out_word = 8'hC0;
		16'h78EA: out_word = 8'hB1;
		16'h78EB: out_word = 8'h0E;
		16'h78EC: out_word = 8'hFD;
		16'h78ED: out_word = 8'hED;
		16'h78EE: out_word = 8'h79;
		16'h78EF: out_word = 8'h7A;
		16'h78F0: out_word = 8'h07;
		16'h78F1: out_word = 8'h07;
		16'h78F2: out_word = 8'h07;
		16'h78F3: out_word = 8'h07;
		16'h78F4: out_word = 8'hE6;
		16'h78F5: out_word = 8'h30;
		16'h78F6: out_word = 8'h83;
		16'h78F7: out_word = 8'hF6;
		16'h78F8: out_word = 8'hC0;
		16'h78F9: out_word = 8'h57;
		16'h78FA: out_word = 8'h1E;
		16'h78FB: out_word = 8'h00;
		16'h78FC: out_word = 8'h3A;
		16'h78FD: out_word = 8'hCE;
		16'h78FE: out_word = 8'h5C;
		16'h78FF: out_word = 8'hA7;
		16'h7900: out_word = 8'h20;
		16'h7901: out_word = 8'h01;
		16'h7902: out_word = 8'hEB;
		16'h7903: out_word = 8'h01;
		16'h7904: out_word = 8'h00;
		16'h7905: out_word = 8'h01;
		16'h7906: out_word = 8'hED;
		16'h7907: out_word = 8'hB0;
		16'h7908: out_word = 8'h3A;
		16'h7909: out_word = 8'h5C;
		16'h790A: out_word = 8'h5B;
		16'h790B: out_word = 8'h01;
		16'h790C: out_word = 8'hFD;
		16'h790D: out_word = 8'h7F;
		16'h790E: out_word = 8'hED;
		16'h790F: out_word = 8'h79;
		16'h7910: out_word = 8'hFB;
		16'h7911: out_word = 8'hC9;
		16'h7912: out_word = 8'h32;
		16'h7913: out_word = 8'hF6;
		16'h7914: out_word = 8'h5C;
		16'h7915: out_word = 8'hFE;
		16'h7916: out_word = 8'h03;
		16'h7917: out_word = 8'hC2;
		16'h7918: out_word = 8'hCE;
		16'h7919: out_word = 8'h3D;
		16'h791A: out_word = 8'hCD;
		16'h791B: out_word = 8'h37;
		16'h791C: out_word = 8'h38;
		16'h791D: out_word = 8'hC2;
		16'h791E: out_word = 8'hE1;
		16'h791F: out_word = 8'h3E;
		16'h7920: out_word = 8'hC9;
		16'h7921: out_word = 8'hCD;
		16'h7922: out_word = 8'h57;
		16'h7923: out_word = 8'h1C;
		16'h7924: out_word = 8'h3A;
		16'h7925: out_word = 8'hF6;
		16'h7926: out_word = 8'h5C;
		16'h7927: out_word = 8'hFE;
		16'h7928: out_word = 8'h03;
		16'h7929: out_word = 8'hC0;
		16'h792A: out_word = 8'hF1;
		16'h792B: out_word = 8'hCD;
		16'h792C: out_word = 8'h54;
		16'h792D: out_word = 8'h39;
		16'h792E: out_word = 8'h11;
		16'h792F: out_word = 8'h00;
		16'h7930: out_word = 8'h00;
		16'h7931: out_word = 8'hED;
		16'h7932: out_word = 8'h53;
		16'h7933: out_word = 8'hF4;
		16'h7934: out_word = 8'h5C;
		16'h7935: out_word = 8'h01;
		16'h7936: out_word = 8'h10;
		16'h7937: out_word = 8'h00;
		16'h7938: out_word = 8'hC5;
		16'h7939: out_word = 8'h3E;
		16'h793A: out_word = 8'hFF;
		16'h793B: out_word = 8'h32;
		16'h793C: out_word = 8'hCE;
		16'h793D: out_word = 8'h5C;
		16'h793E: out_word = 8'h21;
		16'h793F: out_word = 8'h25;
		16'h7940: out_word = 8'h5D;
		16'h7941: out_word = 8'h06;
		16'h7942: out_word = 8'h01;
		16'h7943: out_word = 8'hCD;
		16'h7944: out_word = 8'h1D;
		16'h7945: out_word = 8'h38;
		16'h7946: out_word = 8'hC1;
		16'h7947: out_word = 8'h0B;
		16'h7948: out_word = 8'h78;
		16'h7949: out_word = 8'hB1;
		16'h794A: out_word = 8'h20;
		16'h794B: out_word = 8'hEC;
		16'h794C: out_word = 8'h21;
		16'h794D: out_word = 8'hF0;
		16'h794E: out_word = 8'h07;
		16'h794F: out_word = 8'h3E;
		16'h7950: out_word = 8'h16;
		16'h7951: out_word = 8'hC3;
		16'h7952: out_word = 8'h55;
		16'h7953: out_word = 8'h1F;
		16'h7954: out_word = 8'h21;
		16'h7955: out_word = 8'h25;
		16'h7956: out_word = 8'h5D;
		16'h7957: out_word = 8'h11;
		16'h7958: out_word = 8'h26;
		16'h7959: out_word = 8'h5D;
		16'h795A: out_word = 8'h01;
		16'h795B: out_word = 8'hFF;
		16'h795C: out_word = 8'h00;
		16'h795D: out_word = 8'h70;
		16'h795E: out_word = 8'hED;
		16'h795F: out_word = 8'hB0;
		16'h7960: out_word = 8'hC9;
		16'h7961: out_word = 8'hD5;
		16'h7962: out_word = 8'hE5;
		16'h7963: out_word = 8'hED;
		16'h7964: out_word = 8'h5B;
		16'h7965: out_word = 8'h00;
		16'h7966: out_word = 8'hC0;
		16'h7967: out_word = 8'h2A;
		16'h7968: out_word = 8'hFD;
		16'h7969: out_word = 8'hFF;
		16'h796A: out_word = 8'hE5;
		16'h796B: out_word = 8'h01;
		16'h796C: out_word = 8'hFD;
		16'h796D: out_word = 8'h7F;
		16'h796E: out_word = 8'hED;
		16'h796F: out_word = 8'h43;
		16'h7970: out_word = 8'h00;
		16'h7971: out_word = 8'hC0;
		16'h7972: out_word = 8'hED;
		16'h7973: out_word = 8'h43;
		16'h7974: out_word = 8'hFD;
		16'h7975: out_word = 8'hFF;
		16'h7976: out_word = 8'hAF;
		16'h7977: out_word = 8'hE6;
		16'h7978: out_word = 8'hC7;
		16'h7979: out_word = 8'h3D;
		16'h797A: out_word = 8'hE6;
		16'h797B: out_word = 8'hC7;
		16'h797C: out_word = 8'hF6;
		16'h797D: out_word = 8'h10;
		16'h797E: out_word = 8'hED;
		16'h797F: out_word = 8'h79;
		16'h7980: out_word = 8'h2A;
		16'h7981: out_word = 8'h00;
		16'h7982: out_word = 8'hC0;
		16'h7983: out_word = 8'hED;
		16'h7984: out_word = 8'h42;
		16'h7985: out_word = 8'h20;
		16'h7986: out_word = 8'hF0;
		16'h7987: out_word = 8'h2A;
		16'h7988: out_word = 8'hFD;
		16'h7989: out_word = 8'hFF;
		16'h798A: out_word = 8'hED;
		16'h798B: out_word = 8'h42;
		16'h798C: out_word = 8'h20;
		16'h798D: out_word = 8'hE9;
		16'h798E: out_word = 8'hED;
		16'h798F: out_word = 8'h53;
		16'h7990: out_word = 8'h00;
		16'h7991: out_word = 8'hC0;
		16'h7992: out_word = 8'hE1;
		16'h7993: out_word = 8'h22;
		16'h7994: out_word = 8'hFD;
		16'h7995: out_word = 8'hFF;
		16'h7996: out_word = 8'h32;
		16'h7997: out_word = 8'h5C;
		16'h7998: out_word = 8'h5B;
		16'h7999: out_word = 8'hE1;
		16'h799A: out_word = 8'hD1;
		16'h799B: out_word = 8'hC9;
		16'h799C: out_word = 8'h21;
		16'h799D: out_word = 8'h83;
		16'h799E: out_word = 8'h83;
		16'h799F: out_word = 8'h22;
		16'h79A0: out_word = 8'hC8;
		16'h79A1: out_word = 8'h5C;
		16'h79A2: out_word = 8'h22;
		16'h79A3: out_word = 8'hCA;
		16'h79A4: out_word = 8'h5C;
		16'h79A5: out_word = 8'h3E;
		16'h79A6: out_word = 8'hF7;
		16'h79A7: out_word = 8'hDB;
		16'h79A8: out_word = 8'hFE;
		16'h79A9: out_word = 8'h06;
		16'h79AA: out_word = 8'h00;
		16'h79AB: out_word = 8'h1F;
		16'h79AC: out_word = 8'h30;
		16'h79AD: out_word = 8'h0E;
		16'h79AE: out_word = 8'h04;
		16'h79AF: out_word = 8'h1F;
		16'h79B0: out_word = 8'h30;
		16'h79B1: out_word = 8'h0A;
		16'h79B2: out_word = 8'h04;
		16'h79B3: out_word = 8'h1F;
		16'h79B4: out_word = 8'h30;
		16'h79B5: out_word = 8'h06;
		16'h79B6: out_word = 8'h04;
		16'h79B7: out_word = 8'h1F;
		16'h79B8: out_word = 8'h30;
		16'h79B9: out_word = 8'h02;
		16'h79BA: out_word = 8'h18;
		16'h79BB: out_word = 8'h0E;
		16'h79BC: out_word = 8'h78;
		16'h79BD: out_word = 8'h32;
		16'h79BE: out_word = 8'hF6;
		16'h79BF: out_word = 8'h5C;
		16'h79C0: out_word = 8'h32;
		16'h79C1: out_word = 8'h19;
		16'h79C2: out_word = 8'h5D;
		16'h79C3: out_word = 8'hF6;
		16'h79C4: out_word = 8'h3C;
		16'h79C5: out_word = 8'h32;
		16'h79C6: out_word = 8'h16;
		16'h79C7: out_word = 8'h5D;
		16'h79C8: out_word = 8'hD3;
		16'h79C9: out_word = 8'hFF;
		16'h79CA: out_word = 8'hC3;
		16'h79CB: out_word = 8'h6E;
		16'h79CC: out_word = 8'h10;
		16'h79CD: out_word = 8'hFF;
		16'h79CE: out_word = 8'hFF;
		16'h79CF: out_word = 8'hFF;
		16'h79D0: out_word = 8'hFF;
		16'h79D1: out_word = 8'hFF;
		16'h79D2: out_word = 8'hFF;
		16'h79D3: out_word = 8'hFF;
		16'h79D4: out_word = 8'hFF;
		16'h79D5: out_word = 8'hFF;
		16'h79D6: out_word = 8'hFF;
		16'h79D7: out_word = 8'hFF;
		16'h79D8: out_word = 8'hFF;
		16'h79D9: out_word = 8'hFF;
		16'h79DA: out_word = 8'hFF;
		16'h79DB: out_word = 8'hFF;
		16'h79DC: out_word = 8'hFF;
		16'h79DD: out_word = 8'hFF;
		16'h79DE: out_word = 8'hFF;
		16'h79DF: out_word = 8'hFF;
		16'h79E0: out_word = 8'hFF;
		16'h79E1: out_word = 8'hFF;
		16'h79E2: out_word = 8'hFF;
		16'h79E3: out_word = 8'hFF;
		16'h79E4: out_word = 8'hFF;
		16'h79E5: out_word = 8'hFF;
		16'h79E6: out_word = 8'hFF;
		16'h79E7: out_word = 8'hFF;
		16'h79E8: out_word = 8'hFF;
		16'h79E9: out_word = 8'hFF;
		16'h79EA: out_word = 8'hFF;
		16'h79EB: out_word = 8'hFF;
		16'h79EC: out_word = 8'hFF;
		16'h79ED: out_word = 8'hFF;
		16'h79EE: out_word = 8'hFF;
		16'h79EF: out_word = 8'hFF;
		16'h79F0: out_word = 8'hFF;
		16'h79F1: out_word = 8'hFF;
		16'h79F2: out_word = 8'hFF;
		16'h79F3: out_word = 8'hFF;
		16'h79F4: out_word = 8'hFF;
		16'h79F5: out_word = 8'hFF;
		16'h79F6: out_word = 8'hFF;
		16'h79F7: out_word = 8'hFF;
		16'h79F8: out_word = 8'hFF;
		16'h79F9: out_word = 8'hFF;
		16'h79FA: out_word = 8'hFF;
		16'h79FB: out_word = 8'hFF;
		16'h79FC: out_word = 8'hFF;
		16'h79FD: out_word = 8'hFF;
		16'h79FE: out_word = 8'hFF;
		16'h79FF: out_word = 8'hFF;
		16'h7A00: out_word = 8'hFF;
		16'h7A01: out_word = 8'hFF;
		16'h7A02: out_word = 8'hFF;
		16'h7A03: out_word = 8'hFF;
		16'h7A04: out_word = 8'hFF;
		16'h7A05: out_word = 8'hFF;
		16'h7A06: out_word = 8'hFF;
		16'h7A07: out_word = 8'hFF;
		16'h7A08: out_word = 8'hFF;
		16'h7A09: out_word = 8'hFF;
		16'h7A0A: out_word = 8'hFF;
		16'h7A0B: out_word = 8'hFF;
		16'h7A0C: out_word = 8'hFF;
		16'h7A0D: out_word = 8'hFF;
		16'h7A0E: out_word = 8'hFF;
		16'h7A0F: out_word = 8'hFF;
		16'h7A10: out_word = 8'hFF;
		16'h7A11: out_word = 8'hFF;
		16'h7A12: out_word = 8'hFF;
		16'h7A13: out_word = 8'hFF;
		16'h7A14: out_word = 8'hFF;
		16'h7A15: out_word = 8'hFF;
		16'h7A16: out_word = 8'hFF;
		16'h7A17: out_word = 8'hFF;
		16'h7A18: out_word = 8'hFF;
		16'h7A19: out_word = 8'hFF;
		16'h7A1A: out_word = 8'hFF;
		16'h7A1B: out_word = 8'hFF;
		16'h7A1C: out_word = 8'hFF;
		16'h7A1D: out_word = 8'hFF;
		16'h7A1E: out_word = 8'hFF;
		16'h7A1F: out_word = 8'hFF;
		16'h7A20: out_word = 8'hFF;
		16'h7A21: out_word = 8'hFF;
		16'h7A22: out_word = 8'hFF;
		16'h7A23: out_word = 8'hFF;
		16'h7A24: out_word = 8'hFF;
		16'h7A25: out_word = 8'hFF;
		16'h7A26: out_word = 8'hFF;
		16'h7A27: out_word = 8'hFF;
		16'h7A28: out_word = 8'hFF;
		16'h7A29: out_word = 8'hFF;
		16'h7A2A: out_word = 8'hFF;
		16'h7A2B: out_word = 8'hFF;
		16'h7A2C: out_word = 8'hFF;
		16'h7A2D: out_word = 8'hFF;
		16'h7A2E: out_word = 8'hFF;
		16'h7A2F: out_word = 8'hFF;
		16'h7A30: out_word = 8'hFF;
		16'h7A31: out_word = 8'hFF;
		16'h7A32: out_word = 8'hFF;
		16'h7A33: out_word = 8'hFF;
		16'h7A34: out_word = 8'hFF;
		16'h7A35: out_word = 8'hFF;
		16'h7A36: out_word = 8'hFF;
		16'h7A37: out_word = 8'hFF;
		16'h7A38: out_word = 8'hFF;
		16'h7A39: out_word = 8'hFF;
		16'h7A3A: out_word = 8'hFF;
		16'h7A3B: out_word = 8'hFF;
		16'h7A3C: out_word = 8'hFF;
		16'h7A3D: out_word = 8'hFF;
		16'h7A3E: out_word = 8'hFF;
		16'h7A3F: out_word = 8'hFF;
		16'h7A40: out_word = 8'hFF;
		16'h7A41: out_word = 8'hFF;
		16'h7A42: out_word = 8'hFF;
		16'h7A43: out_word = 8'hFF;
		16'h7A44: out_word = 8'hFF;
		16'h7A45: out_word = 8'hFF;
		16'h7A46: out_word = 8'hFF;
		16'h7A47: out_word = 8'hFF;
		16'h7A48: out_word = 8'hFF;
		16'h7A49: out_word = 8'hFF;
		16'h7A4A: out_word = 8'hFF;
		16'h7A4B: out_word = 8'hFF;
		16'h7A4C: out_word = 8'hFF;
		16'h7A4D: out_word = 8'hFF;
		16'h7A4E: out_word = 8'hFF;
		16'h7A4F: out_word = 8'hFF;
		16'h7A50: out_word = 8'hFF;
		16'h7A51: out_word = 8'hFF;
		16'h7A52: out_word = 8'hFF;
		16'h7A53: out_word = 8'hFF;
		16'h7A54: out_word = 8'hFF;
		16'h7A55: out_word = 8'hFF;
		16'h7A56: out_word = 8'hFF;
		16'h7A57: out_word = 8'hFF;
		16'h7A58: out_word = 8'hFF;
		16'h7A59: out_word = 8'hFF;
		16'h7A5A: out_word = 8'hFF;
		16'h7A5B: out_word = 8'hFF;
		16'h7A5C: out_word = 8'hFF;
		16'h7A5D: out_word = 8'hFF;
		16'h7A5E: out_word = 8'hFF;
		16'h7A5F: out_word = 8'hFF;
		16'h7A60: out_word = 8'hFF;
		16'h7A61: out_word = 8'hFF;
		16'h7A62: out_word = 8'hFF;
		16'h7A63: out_word = 8'hFF;
		16'h7A64: out_word = 8'hFF;
		16'h7A65: out_word = 8'hFF;
		16'h7A66: out_word = 8'hFF;
		16'h7A67: out_word = 8'hFF;
		16'h7A68: out_word = 8'hFF;
		16'h7A69: out_word = 8'hFF;
		16'h7A6A: out_word = 8'hFF;
		16'h7A6B: out_word = 8'hFF;
		16'h7A6C: out_word = 8'hFF;
		16'h7A6D: out_word = 8'hFF;
		16'h7A6E: out_word = 8'hFF;
		16'h7A6F: out_word = 8'hFF;
		16'h7A70: out_word = 8'hFF;
		16'h7A71: out_word = 8'hFF;
		16'h7A72: out_word = 8'hFF;
		16'h7A73: out_word = 8'hFF;
		16'h7A74: out_word = 8'hFF;
		16'h7A75: out_word = 8'hFF;
		16'h7A76: out_word = 8'hFF;
		16'h7A77: out_word = 8'hFF;
		16'h7A78: out_word = 8'hFF;
		16'h7A79: out_word = 8'hFF;
		16'h7A7A: out_word = 8'hFF;
		16'h7A7B: out_word = 8'hFF;
		16'h7A7C: out_word = 8'hFF;
		16'h7A7D: out_word = 8'hFF;
		16'h7A7E: out_word = 8'hFF;
		16'h7A7F: out_word = 8'hFF;
		16'h7A80: out_word = 8'hFF;
		16'h7A81: out_word = 8'hFF;
		16'h7A82: out_word = 8'hFF;
		16'h7A83: out_word = 8'hFF;
		16'h7A84: out_word = 8'hFF;
		16'h7A85: out_word = 8'hFF;
		16'h7A86: out_word = 8'hFF;
		16'h7A87: out_word = 8'hFF;
		16'h7A88: out_word = 8'hFF;
		16'h7A89: out_word = 8'hFF;
		16'h7A8A: out_word = 8'hFF;
		16'h7A8B: out_word = 8'hFF;
		16'h7A8C: out_word = 8'hFF;
		16'h7A8D: out_word = 8'hFF;
		16'h7A8E: out_word = 8'hFF;
		16'h7A8F: out_word = 8'hFF;
		16'h7A90: out_word = 8'hFF;
		16'h7A91: out_word = 8'hFF;
		16'h7A92: out_word = 8'hFF;
		16'h7A93: out_word = 8'hFF;
		16'h7A94: out_word = 8'hFF;
		16'h7A95: out_word = 8'hFF;
		16'h7A96: out_word = 8'hFF;
		16'h7A97: out_word = 8'hFF;
		16'h7A98: out_word = 8'hFF;
		16'h7A99: out_word = 8'hFF;
		16'h7A9A: out_word = 8'hFF;
		16'h7A9B: out_word = 8'hFF;
		16'h7A9C: out_word = 8'hFF;
		16'h7A9D: out_word = 8'hFF;
		16'h7A9E: out_word = 8'hFF;
		16'h7A9F: out_word = 8'hFF;
		16'h7AA0: out_word = 8'hFF;
		16'h7AA1: out_word = 8'hFF;
		16'h7AA2: out_word = 8'hFF;
		16'h7AA3: out_word = 8'hFF;
		16'h7AA4: out_word = 8'hFF;
		16'h7AA5: out_word = 8'hFF;
		16'h7AA6: out_word = 8'hFF;
		16'h7AA7: out_word = 8'hFF;
		16'h7AA8: out_word = 8'hFF;
		16'h7AA9: out_word = 8'hFF;
		16'h7AAA: out_word = 8'hFF;
		16'h7AAB: out_word = 8'hFF;
		16'h7AAC: out_word = 8'hFF;
		16'h7AAD: out_word = 8'hFF;
		16'h7AAE: out_word = 8'hFF;
		16'h7AAF: out_word = 8'hFF;
		16'h7AB0: out_word = 8'hFF;
		16'h7AB1: out_word = 8'hFF;
		16'h7AB2: out_word = 8'hFF;
		16'h7AB3: out_word = 8'hFF;
		16'h7AB4: out_word = 8'hFF;
		16'h7AB5: out_word = 8'hFF;
		16'h7AB6: out_word = 8'hFF;
		16'h7AB7: out_word = 8'hFF;
		16'h7AB8: out_word = 8'hFF;
		16'h7AB9: out_word = 8'hFF;
		16'h7ABA: out_word = 8'hFF;
		16'h7ABB: out_word = 8'hFF;
		16'h7ABC: out_word = 8'hFF;
		16'h7ABD: out_word = 8'hFF;
		16'h7ABE: out_word = 8'hFF;
		16'h7ABF: out_word = 8'hFF;
		16'h7AC0: out_word = 8'hFF;
		16'h7AC1: out_word = 8'hFF;
		16'h7AC2: out_word = 8'hFF;
		16'h7AC3: out_word = 8'hFF;
		16'h7AC4: out_word = 8'hFF;
		16'h7AC5: out_word = 8'hFF;
		16'h7AC6: out_word = 8'hFF;
		16'h7AC7: out_word = 8'hFF;
		16'h7AC8: out_word = 8'hFF;
		16'h7AC9: out_word = 8'hFF;
		16'h7ACA: out_word = 8'hFF;
		16'h7ACB: out_word = 8'hFF;
		16'h7ACC: out_word = 8'hFF;
		16'h7ACD: out_word = 8'hFF;
		16'h7ACE: out_word = 8'hFF;
		16'h7ACF: out_word = 8'hFF;
		16'h7AD0: out_word = 8'hFF;
		16'h7AD1: out_word = 8'hFF;
		16'h7AD2: out_word = 8'hFF;
		16'h7AD3: out_word = 8'hFF;
		16'h7AD4: out_word = 8'hFF;
		16'h7AD5: out_word = 8'hFF;
		16'h7AD6: out_word = 8'hFF;
		16'h7AD7: out_word = 8'hFF;
		16'h7AD8: out_word = 8'hFF;
		16'h7AD9: out_word = 8'hFF;
		16'h7ADA: out_word = 8'hFF;
		16'h7ADB: out_word = 8'h01;
		16'h7ADC: out_word = 8'hFF;
		16'h7ADD: out_word = 8'hF4;
		16'h7ADE: out_word = 8'hE7;
		16'h7ADF: out_word = 8'hAF;
		16'h7AE0: out_word = 8'h1E;
		16'h7AE1: out_word = 8'h3E;
		16'h7AE2: out_word = 8'h01;
		16'h7AE3: out_word = 8'hE7;
		16'h7AE4: out_word = 8'h9B;
		16'h7AE5: out_word = 8'h22;
		16'h7AE6: out_word = 8'hF3;
		16'h7AE7: out_word = 8'h21;
		16'h7AE8: out_word = 8'h00;
		16'h7AE9: out_word = 8'h0E;
		16'h7AEA: out_word = 8'h11;
		16'h7AEB: out_word = 8'h00;
		16'h7AEC: out_word = 8'hF5;
		16'h7AED: out_word = 8'h01;
		16'h7AEE: out_word = 8'hF5;
		16'h7AEF: out_word = 8'h01;
		16'h7AF0: out_word = 8'hD5;
		16'h7AF1: out_word = 8'hED;
		16'h7AF2: out_word = 8'hB0;
		16'h7AF3: out_word = 8'h21;
		16'h7AF4: out_word = 8'h4D;
		16'h7AF5: out_word = 8'h34;
		16'h7AF6: out_word = 8'h01;
		16'h7AF7: out_word = 8'h34;
		16'h7AF8: out_word = 8'h03;
		16'h7AF9: out_word = 8'hED;
		16'h7AFA: out_word = 8'hB0;
		16'h7AFB: out_word = 8'hFD;
		16'h7AFC: out_word = 8'hCB;
		16'h7AFD: out_word = 8'h01;
		16'h7AFE: out_word = 8'hDE;
		16'h7AFF: out_word = 8'hC9;
		16'h7B00: out_word = 8'h2A;
		16'h7B01: out_word = 8'hE1;
		16'h7B02: out_word = 8'h5C;
		16'h7B03: out_word = 8'h7E;
		16'h7B04: out_word = 8'hFE;
		16'h7B05: out_word = 8'h00;
		16'h7B06: out_word = 8'hC8;
		16'h7B07: out_word = 8'hFE;
		16'h7B08: out_word = 8'h01;
		16'h7B09: out_word = 8'h28;
		16'h7B0A: out_word = 8'h03;
		16'h7B0B: out_word = 8'hCD;
		16'h7B0C: out_word = 8'h14;
		16'h7B0D: out_word = 8'h3B;
		16'h7B0E: out_word = 8'h11;
		16'h7B0F: out_word = 8'h10;
		16'h7B10: out_word = 8'h00;
		16'h7B11: out_word = 8'h19;
		16'h7B12: out_word = 8'h18;
		16'h7B13: out_word = 8'hEF;
		16'h7B14: out_word = 8'hE5;
		16'h7B15: out_word = 8'h11;
		16'h7B16: out_word = 8'h0D;
		16'h7B17: out_word = 8'h00;
		16'h7B18: out_word = 8'h19;
		16'h7B19: out_word = 8'h4E;
		16'h7B1A: out_word = 8'h23;
		16'h7B1B: out_word = 8'h5E;
		16'h7B1C: out_word = 8'h23;
		16'h7B1D: out_word = 8'h56;
		16'h7B1E: out_word = 8'h2A;
		16'h7B1F: out_word = 8'hD7;
		16'h7B20: out_word = 8'h5C;
		16'h7B21: out_word = 8'hA7;
		16'h7B22: out_word = 8'hED;
		16'h7B23: out_word = 8'h52;
		16'h7B24: out_word = 8'h19;
		16'h7B25: out_word = 8'h28;
		16'h7B26: out_word = 8'h2F;
		16'h7B27: out_word = 8'hED;
		16'h7B28: out_word = 8'h53;
		16'h7B29: out_word = 8'hD5;
		16'h7B2A: out_word = 8'h5C;
		16'h7B2B: out_word = 8'h79;
		16'h7B2C: out_word = 8'h32;
		16'h7B2D: out_word = 8'hD3;
		16'h7B2E: out_word = 8'h5C;
		16'h7B2F: out_word = 8'hCD;
		16'h7B30: out_word = 8'hA5;
		16'h7B31: out_word = 8'h17;
		16'h7B32: out_word = 8'hE1;
		16'h7B33: out_word = 8'hE5;
		16'h7B34: out_word = 8'hED;
		16'h7B35: out_word = 8'h5B;
		16'h7B36: out_word = 8'hDF;
		16'h7B37: out_word = 8'h5C;
		16'h7B38: out_word = 8'h01;
		16'h7B39: out_word = 8'h10;
		16'h7B3A: out_word = 8'h00;
		16'h7B3B: out_word = 8'hED;
		16'h7B3C: out_word = 8'hB0;
		16'h7B3D: out_word = 8'hED;
		16'h7B3E: out_word = 8'h53;
		16'h7B3F: out_word = 8'hDF;
		16'h7B40: out_word = 8'h5C;
		16'h7B41: out_word = 8'hEB;
		16'h7B42: out_word = 8'hED;
		16'h7B43: out_word = 8'h5B;
		16'h7B44: out_word = 8'hDD;
		16'h7B45: out_word = 8'h5C;
		16'h7B46: out_word = 8'h2B;
		16'h7B47: out_word = 8'h72;
		16'h7B48: out_word = 8'h2B;
		16'h7B49: out_word = 8'h73;
		16'h7B4A: out_word = 8'h2A;
		16'h7B4B: out_word = 8'hD7;
		16'h7B4C: out_word = 8'h5C;
		16'h7B4D: out_word = 8'h22;
		16'h7B4E: out_word = 8'hDD;
		16'h7B4F: out_word = 8'h5C;
		16'h7B50: out_word = 8'h21;
		16'h7B51: out_word = 8'hE3;
		16'h7B52: out_word = 8'h5C;
		16'h7B53: out_word = 8'h34;
		16'h7B54: out_word = 8'hE1;
		16'h7B55: out_word = 8'hC9;
		16'h7B56: out_word = 8'h79;
		16'h7B57: out_word = 8'hE6;
		16'h7B58: out_word = 8'h0F;
		16'h7B59: out_word = 8'h83;
		16'h7B5A: out_word = 8'hCB;
		16'h7B5B: out_word = 8'h67;
		16'h7B5C: out_word = 8'hCB;
		16'h7B5D: out_word = 8'hA7;
		16'h7B5E: out_word = 8'h5F;
		16'h7B5F: out_word = 8'h28;
		16'h7B60: out_word = 8'h01;
		16'h7B61: out_word = 8'h14;
		16'h7B62: out_word = 8'h79;
		16'h7B63: out_word = 8'hCB;
		16'h7B64: out_word = 8'h0F;
		16'h7B65: out_word = 8'hCB;
		16'h7B66: out_word = 8'h0F;
		16'h7B67: out_word = 8'hCB;
		16'h7B68: out_word = 8'h0F;
		16'h7B69: out_word = 8'hCB;
		16'h7B6A: out_word = 8'h0F;
		16'h7B6B: out_word = 8'hE6;
		16'h7B6C: out_word = 8'h0F;
		16'h7B6D: out_word = 8'h82;
		16'h7B6E: out_word = 8'h57;
		16'h7B6F: out_word = 8'hED;
		16'h7B70: out_word = 8'h53;
		16'h7B71: out_word = 8'hD7;
		16'h7B72: out_word = 8'h5C;
		16'h7B73: out_word = 8'h18;
		16'h7B74: out_word = 8'hBD;
		16'h7B75: out_word = 8'hFF;
		16'h7B76: out_word = 8'hFF;
		16'h7B77: out_word = 8'hFF;
		16'h7B78: out_word = 8'hFF;
		16'h7B79: out_word = 8'hFF;
		16'h7B7A: out_word = 8'hFF;
		16'h7B7B: out_word = 8'hFF;
		16'h7B7C: out_word = 8'hFF;
		16'h7B7D: out_word = 8'hFF;
		16'h7B7E: out_word = 8'hFF;
		16'h7B7F: out_word = 8'hFF;
		16'h7B80: out_word = 8'hFD;
		16'h7B81: out_word = 8'hCB;
		16'h7B82: out_word = 8'h01;
		16'h7B83: out_word = 8'hAE;
		16'h7B84: out_word = 8'hE7;
		16'h7B85: out_word = 8'hD4;
		16'h7B86: out_word = 8'h15;
		16'h7B87: out_word = 8'hFE;
		16'h7B88: out_word = 8'h07;
		16'h7B89: out_word = 8'h20;
		16'h7B8A: out_word = 8'h22;
		16'h7B8B: out_word = 8'h21;
		16'h7B8C: out_word = 8'hC8;
		16'h7B8D: out_word = 8'h00;
		16'h7B8E: out_word = 8'h54;
		16'h7B8F: out_word = 8'hFD;
		16'h7B90: out_word = 8'h5E;
		16'h7B91: out_word = 8'hFF;
		16'h7B92: out_word = 8'hE7;
		16'h7B93: out_word = 8'hB5;
		16'h7B94: out_word = 8'h03;
		16'h7B95: out_word = 8'hCD;
		16'h7B96: out_word = 8'h2A;
		16'h7B97: out_word = 8'h21;
		16'h7B98: out_word = 8'h2A;
		16'h7B99: out_word = 8'h59;
		16'h7B9A: out_word = 8'h5C;
		16'h7B9B: out_word = 8'h3E;
		16'h7B9C: out_word = 8'h0D;
		16'h7B9D: out_word = 8'h01;
		16'h7B9E: out_word = 8'h00;
		16'h7B9F: out_word = 8'h00;
		16'h7BA0: out_word = 8'hED;
		16'h7BA1: out_word = 8'hB1;
		16'h7BA2: out_word = 8'h2B;
		16'h7BA3: out_word = 8'h22;
		16'h7BA4: out_word = 8'h5B;
		16'h7BA5: out_word = 8'h5C;
		16'h7BA6: out_word = 8'h23;
		16'h7BA7: out_word = 8'h23;
		16'h7BA8: out_word = 8'h36;
		16'h7BA9: out_word = 8'h80;
		16'h7BAA: out_word = 8'hE7;
		16'h7BAB: out_word = 8'hD4;
		16'h7BAC: out_word = 8'h15;
		16'h7BAD: out_word = 8'hF5;
		16'h7BAE: out_word = 8'h21;
		16'h7BAF: out_word = 8'hC8;
		16'h7BB0: out_word = 8'h00;
		16'h7BB1: out_word = 8'h54;
		16'h7BB2: out_word = 8'hFD;
		16'h7BB3: out_word = 8'h5E;
		16'h7BB4: out_word = 8'hFF;
		16'h7BB5: out_word = 8'hE7;
		16'h7BB6: out_word = 8'hB5;
		16'h7BB7: out_word = 8'h03;
		16'h7BB8: out_word = 8'hF1;
		16'h7BB9: out_word = 8'hFE;
		16'h7BBA: out_word = 8'h18;
		16'h7BBB: out_word = 8'h30;
		16'h7BBC: out_word = 8'h0D;
		16'h7BBD: out_word = 8'hFE;
		16'h7BBE: out_word = 8'h07;
		16'h7BBF: out_word = 8'h38;
		16'h7BC0: out_word = 8'h09;
		16'h7BC1: out_word = 8'hFE;
		16'h7BC2: out_word = 8'h10;
		16'h7BC3: out_word = 8'h38;
		16'h7BC4: out_word = 8'h0A;
		16'h7BC5: out_word = 8'hE7;
		16'h7BC6: out_word = 8'h58;
		16'h7BC7: out_word = 8'h0F;
		16'h7BC8: out_word = 8'h18;
		16'h7BC9: out_word = 8'hE0;
		16'h7BCA: out_word = 8'hE7;
		16'h7BCB: out_word = 8'h81;
		16'h7BCC: out_word = 8'h0F;
		16'h7BCD: out_word = 8'h18;
		16'h7BCE: out_word = 8'hDB;
		16'h7BCF: out_word = 8'hFE;
		16'h7BD0: out_word = 8'h07;
		16'h7BD1: out_word = 8'h28;
		16'h7BD2: out_word = 8'hD7;
		16'h7BD3: out_word = 8'hFE;
		16'h7BD4: out_word = 8'h0D;
		16'h7BD5: out_word = 8'hC8;
		16'h7BD6: out_word = 8'hFE;
		16'h7BD7: out_word = 8'h0A;
		16'h7BD8: out_word = 8'h28;
		16'h7BD9: out_word = 8'hD0;
		16'h7BDA: out_word = 8'hFE;
		16'h7BDB: out_word = 8'h0B;
		16'h7BDC: out_word = 8'h28;
		16'h7BDD: out_word = 8'hCC;
		16'h7BDE: out_word = 8'hE7;
		16'h7BDF: out_word = 8'h92;
		16'h7BE0: out_word = 8'h0F;
		16'h7BE1: out_word = 8'h18;
		16'h7BE2: out_word = 8'hC7;
		16'h7BE3: out_word = 8'hFF;
		16'h7BE4: out_word = 8'hFF;
		16'h7BE5: out_word = 8'hFF;
		16'h7BE6: out_word = 8'hFF;
		16'h7BE7: out_word = 8'hFF;
		16'h7BE8: out_word = 8'hFF;
		16'h7BE9: out_word = 8'hFF;
		16'h7BEA: out_word = 8'hFF;
		16'h7BEB: out_word = 8'hFF;
		16'h7BEC: out_word = 8'hFF;
		16'h7BED: out_word = 8'hFF;
		16'h7BEE: out_word = 8'hFF;
		16'h7BEF: out_word = 8'hFF;
		16'h7BF0: out_word = 8'hCD;
		16'h7BF1: out_word = 8'h9F;
		16'h7BF2: out_word = 8'h1D;
		16'h7BF3: out_word = 8'hC3;
		16'h7BF4: out_word = 8'h39;
		16'h7BF5: out_word = 8'h02;
		16'h7BF6: out_word = 8'h21;
		16'h7BF7: out_word = 8'h06;
		16'h7BF8: out_word = 8'h5E;
		16'h7BF9: out_word = 8'h3E;
		16'h7BFA: out_word = 8'hFF;
		16'h7BFB: out_word = 8'h32;
		16'h7BFC: out_word = 8'h0E;
		16'h7BFD: out_word = 8'h5D;
		16'h7BFE: out_word = 8'hC9;
		16'h7BFF: out_word = 8'hFF;
		16'h7C00: out_word = 8'hFF;
		16'h7C01: out_word = 8'h18;
		16'h7C02: out_word = 8'h03;
		16'h7C03: out_word = 8'hFF;
		16'h7C04: out_word = 8'h18;
		16'h7C05: out_word = 8'h03;
		16'h7C06: out_word = 8'hC3;
		16'h7C07: out_word = 8'h00;
		16'h7C08: out_word = 8'h3D;
		16'h7C09: out_word = 8'hC3;
		16'h7C0A: out_word = 8'h03;
		16'h7C0B: out_word = 8'h3D;
		16'h7C0C: out_word = 8'hFF;
		16'h7C0D: out_word = 8'hFF;
		16'h7C0E: out_word = 8'hFF;
		16'h7C0F: out_word = 8'hFF;
		16'h7C10: out_word = 8'h4A;
		16'h7C11: out_word = 8'hED;
		16'h7C12: out_word = 8'h59;
		16'h7C13: out_word = 8'hC9;
		16'h7C14: out_word = 8'h4A;
		16'h7C15: out_word = 8'hED;
		16'h7C16: out_word = 8'h58;
		16'h7C17: out_word = 8'hC9;
		16'h7C18: out_word = 8'h0E;
		16'h7C19: out_word = 8'h7F;
		16'h7C1A: out_word = 8'hC3;
		16'h7C1B: out_word = 8'hBA;
		16'h7C1C: out_word = 8'h3F;
		16'h7C1D: out_word = 8'h0E;
		16'h7C1E: out_word = 8'h7F;
		16'h7C1F: out_word = 8'hC3;
		16'h7C20: out_word = 8'hD5;
		16'h7C21: out_word = 8'h3F;
		16'h7C22: out_word = 8'hFF;
		16'h7C23: out_word = 8'hFF;
		16'h7C24: out_word = 8'hFF;
		16'h7C25: out_word = 8'hFF;
		16'h7C26: out_word = 8'hFF;
		16'h7C27: out_word = 8'hFF;
		16'h7C28: out_word = 8'hFF;
		16'h7C29: out_word = 8'hFF;
		16'h7C2A: out_word = 8'hFF;
		16'h7C2B: out_word = 8'hFF;
		16'h7C2C: out_word = 8'hFF;
		16'h7C2D: out_word = 8'hFF;
		16'h7C2E: out_word = 8'hFF;
		16'h7C2F: out_word = 8'hFF;
		16'h7C30: out_word = 8'hDB;
		16'h7C31: out_word = 8'h1F;
		16'h7C32: out_word = 8'hC9;
		16'h7C33: out_word = 8'hFF;
		16'h7C34: out_word = 8'hFF;
		16'h7C35: out_word = 8'hFF;
		16'h7C36: out_word = 8'hFF;
		16'h7C37: out_word = 8'hFF;
		16'h7C38: out_word = 8'hFF;
		16'h7C39: out_word = 8'hFF;
		16'h7C3A: out_word = 8'hFF;
		16'h7C3B: out_word = 8'hFF;
		16'h7C3C: out_word = 8'hFF;
		16'h7C3D: out_word = 8'hFF;
		16'h7C3E: out_word = 8'hFF;
		16'h7C3F: out_word = 8'hFF;
		16'h7C40: out_word = 8'hFF;
		16'h7C41: out_word = 8'hFF;
		16'h7C42: out_word = 8'hFF;
		16'h7C43: out_word = 8'hFF;
		16'h7C44: out_word = 8'hFF;
		16'h7C45: out_word = 8'hFF;
		16'h7C46: out_word = 8'hFF;
		16'h7C47: out_word = 8'hFF;
		16'h7C48: out_word = 8'hC3;
		16'h7C49: out_word = 8'h9A;
		16'h7C4A: out_word = 8'h37;
		16'h7C4B: out_word = 8'h3E;
		16'h7C4C: out_word = 8'h07;
		16'h7C4D: out_word = 8'hC3;
		16'h7C4E: out_word = 8'h09;
		16'h7C4F: out_word = 8'h00;
		16'h7C50: out_word = 8'h31;
		16'h7C51: out_word = 8'hFF;
		16'h7C52: out_word = 8'h5B;
		16'h7C53: out_word = 8'h3E;
		16'h7C54: out_word = 8'h1F;
		16'h7C55: out_word = 8'hCD;
		16'h7C56: out_word = 8'hC5;
		16'h7C57: out_word = 8'h3C;
		16'h7C58: out_word = 8'h21;
		16'h7C59: out_word = 8'h00;
		16'h7C5A: out_word = 8'hC0;
		16'h7C5B: out_word = 8'h7E;
		16'h7C5C: out_word = 8'hFE;
		16'h7C5D: out_word = 8'hC3;
		16'h7C5E: out_word = 8'h20;
		16'h7C5F: out_word = 8'hE8;
		16'h7C60: out_word = 8'hAF;
		16'h7C61: out_word = 8'h86;
		16'h7C62: out_word = 8'hCE;
		16'h7C63: out_word = 8'h00;
		16'h7C64: out_word = 8'h23;
		16'h7C65: out_word = 8'hCB;
		16'h7C66: out_word = 8'h7C;
		16'h7C67: out_word = 8'h20;
		16'h7C68: out_word = 8'hF8;
		16'h7C69: out_word = 8'h3D;
		16'h7C6A: out_word = 8'h20;
		16'h7C6B: out_word = 8'hDC;
		16'h7C6C: out_word = 8'h3E;
		16'h7C6D: out_word = 8'hAA;
		16'h7C6E: out_word = 8'h2B;
		16'h7C6F: out_word = 8'hBE;
		16'h7C70: out_word = 8'h20;
		16'h7C71: out_word = 8'hD6;
		16'h7C72: out_word = 8'h2F;
		16'h7C73: out_word = 8'h2B;
		16'h7C74: out_word = 8'hBE;
		16'h7C75: out_word = 8'h20;
		16'h7C76: out_word = 8'hD1;
		16'h7C77: out_word = 8'h21;
		16'h7C78: out_word = 8'h00;
		16'h7C79: out_word = 8'hD0;
		16'h7C7A: out_word = 8'h11;
		16'h7C7B: out_word = 8'h00;
		16'h7C7C: out_word = 8'h5B;
		16'h7C7D: out_word = 8'h01;
		16'h7C7E: out_word = 8'h00;
		16'h7C7F: out_word = 8'h25;
		16'h7C80: out_word = 8'hED;
		16'h7C81: out_word = 8'hB0;
		16'h7C82: out_word = 8'h31;
		16'h7C83: out_word = 8'h00;
		16'h7C84: out_word = 8'h5F;
		16'h7C85: out_word = 8'h3E;
		16'h7C86: out_word = 8'h1E;
		16'h7C87: out_word = 8'hCD;
		16'h7C88: out_word = 8'hC5;
		16'h7C89: out_word = 8'h3C;
		16'h7C8A: out_word = 8'hCD;
		16'h7C8B: out_word = 8'hDF;
		16'h7C8C: out_word = 8'h3C;
		16'h7C8D: out_word = 8'h3E;
		16'h7C8E: out_word = 8'h03;
		16'h7C8F: out_word = 8'hCD;
		16'h7C90: out_word = 8'hC5;
		16'h7C91: out_word = 8'h3C;
		16'h7C92: out_word = 8'hCD;
		16'h7C93: out_word = 8'hDA;
		16'h7C94: out_word = 8'h3C;
		16'h7C95: out_word = 8'h3E;
		16'h7C96: out_word = 8'h1D;
		16'h7C97: out_word = 8'hCD;
		16'h7C98: out_word = 8'hC5;
		16'h7C99: out_word = 8'h3C;
		16'h7C9A: out_word = 8'hCD;
		16'h7C9B: out_word = 8'hDF;
		16'h7C9C: out_word = 8'h3C;
		16'h7C9D: out_word = 8'h3E;
		16'h7C9E: out_word = 8'h01;
		16'h7C9F: out_word = 8'hCD;
		16'h7CA0: out_word = 8'hC5;
		16'h7CA1: out_word = 8'h3C;
		16'h7CA2: out_word = 8'hCD;
		16'h7CA3: out_word = 8'hDA;
		16'h7CA4: out_word = 8'h3C;
		16'h7CA5: out_word = 8'h3E;
		16'h7CA6: out_word = 8'h1C;
		16'h7CA7: out_word = 8'hCD;
		16'h7CA8: out_word = 8'hC5;
		16'h7CA9: out_word = 8'h3C;
		16'h7CAA: out_word = 8'hCD;
		16'h7CAB: out_word = 8'hDF;
		16'h7CAC: out_word = 8'h3C;
		16'h7CAD: out_word = 8'hAF;
		16'h7CAE: out_word = 8'hCD;
		16'h7CAF: out_word = 8'hC5;
		16'h7CB0: out_word = 8'h3C;
		16'h7CB1: out_word = 8'hCD;
		16'h7CB2: out_word = 8'hDA;
		16'h7CB3: out_word = 8'h3C;
		16'h7CB4: out_word = 8'h3E;
		16'h7CB5: out_word = 8'h1B;
		16'h7CB6: out_word = 8'hCD;
		16'h7CB7: out_word = 8'hC5;
		16'h7CB8: out_word = 8'h3C;
		16'h7CB9: out_word = 8'hCD;
		16'h7CBA: out_word = 8'hDF;
		16'h7CBB: out_word = 8'h3C;
		16'h7CBC: out_word = 8'hAF;
		16'h7CBD: out_word = 8'hCD;
		16'h7CBE: out_word = 8'hC5;
		16'h7CBF: out_word = 8'h3C;
		16'h7CC0: out_word = 8'hED;
		16'h7CC1: out_word = 8'h7B;
		16'h7CC2: out_word = 8'h73;
		16'h7CC3: out_word = 8'h5B;
		16'h7CC4: out_word = 8'hC9;
		16'h7CC5: out_word = 8'hF5;
		16'h7CC6: out_word = 8'h17;
		16'h7CC7: out_word = 8'h17;
		16'h7CC8: out_word = 8'h17;
		16'h7CC9: out_word = 8'hE6;
		16'h7CCA: out_word = 8'hC0;
		16'h7CCB: out_word = 8'h4F;
		16'h7CCC: out_word = 8'hF1;
		16'h7CCD: out_word = 8'hE6;
		16'h7CCE: out_word = 8'h27;
		16'h7CCF: out_word = 8'hB1;
		16'h7CD0: out_word = 8'hF6;
		16'h7CD1: out_word = 8'h10;
		16'h7CD2: out_word = 8'h01;
		16'h7CD3: out_word = 8'hFD;
		16'h7CD4: out_word = 8'h7F;
		16'h7CD5: out_word = 8'hED;
		16'h7CD6: out_word = 8'h79;
		16'h7CD7: out_word = 8'hC9;
		16'h7CD8: out_word = 8'hFF;
		16'h7CD9: out_word = 8'hFF;
		16'h7CDA: out_word = 8'h3E;
		16'h7CDB: out_word = 8'hFF;
		16'h7CDC: out_word = 8'hB7;
		16'h7CDD: out_word = 8'h18;
		16'h7CDE: out_word = 8'h01;
		16'h7CDF: out_word = 8'hAF;
		16'h7CE0: out_word = 8'h21;
		16'h7CE1: out_word = 8'h00;
		16'h7CE2: out_word = 8'hC0;
		16'h7CE3: out_word = 8'h11;
		16'h7CE4: out_word = 8'h00;
		16'h7CE5: out_word = 8'h80;
		16'h7CE6: out_word = 8'h01;
		16'h7CE7: out_word = 8'h00;
		16'h7CE8: out_word = 8'h40;
		16'h7CE9: out_word = 8'h28;
		16'h7CEA: out_word = 8'h01;
		16'h7CEB: out_word = 8'hEB;
		16'h7CEC: out_word = 8'hED;
		16'h7CED: out_word = 8'hB0;
		16'h7CEE: out_word = 8'hC9;
		16'h7CEF: out_word = 8'hFF;
		16'h7CF0: out_word = 8'hFF;
		16'h7CF1: out_word = 8'hFF;
		16'h7CF2: out_word = 8'hFF;
		16'h7CF3: out_word = 8'hFF;
		16'h7CF4: out_word = 8'hFF;
		16'h7CF5: out_word = 8'hFF;
		16'h7CF6: out_word = 8'hFF;
		16'h7CF7: out_word = 8'hFF;
		16'h7CF8: out_word = 8'hFF;
		16'h7CF9: out_word = 8'hFF;
		16'h7CFA: out_word = 8'hC3;
		16'h7CFB: out_word = 8'hF1;
		16'h7CFC: out_word = 8'h20;
		16'h7CFD: out_word = 8'hC3;
		16'h7CFE: out_word = 8'h3C;
		16'h7CFF: out_word = 8'h28;
		16'h7D00: out_word = 8'h00;
		16'h7D01: out_word = 8'h18;
		16'h7D02: out_word = 8'h2E;
		16'h7D03: out_word = 8'h00;
		16'h7D04: out_word = 8'h18;
		16'h7D05: out_word = 8'h14;
		16'h7D06: out_word = 8'h00;
		16'h7D07: out_word = 8'hC3;
		16'h7D08: out_word = 8'hEF;
		16'h7D09: out_word = 8'h25;
		16'h7D0A: out_word = 8'hC3;
		16'h7D0B: out_word = 8'h4A;
		16'h7D0C: out_word = 8'h24;
		16'h7D0D: out_word = 8'h00;
		16'h7D0E: out_word = 8'h18;
		16'h7D0F: out_word = 8'hFA;
		16'h7D10: out_word = 8'h00;
		16'h7D11: out_word = 8'h18;
		16'h7D12: out_word = 8'hE7;
		16'h7D13: out_word = 8'h00;
		16'h7D14: out_word = 8'h18;
		16'h7D15: out_word = 8'hE7;
		16'h7D16: out_word = 8'h00;
		16'h7D17: out_word = 8'hC3;
		16'h7D18: out_word = 8'h49;
		16'h7D19: out_word = 8'h34;
		16'h7D1A: out_word = 8'hCD;
		16'h7D1B: out_word = 8'h21;
		16'h7D1C: out_word = 8'h3D;
		16'h7D1D: out_word = 8'hE5;
		16'h7D1E: out_word = 8'hC3;
		16'h7D1F: out_word = 8'h6C;
		16'h7D20: out_word = 8'h01;
		16'h7D21: out_word = 8'hCD;
		16'h7D22: out_word = 8'hF3;
		16'h7D23: out_word = 8'h31;
		16'h7D24: out_word = 8'h00;
		16'h7D25: out_word = 8'h00;
		16'h7D26: out_word = 8'hDC;
		16'h7D27: out_word = 8'h4C;
		16'h7D28: out_word = 8'h3D;
		16'h7D29: out_word = 8'h21;
		16'h7D2A: out_word = 8'hC2;
		16'h7D2B: out_word = 8'h5C;
		16'h7D2C: out_word = 8'hC9;
		16'h7D2D: out_word = 8'h00;
		16'h7D2E: out_word = 8'h00;
		16'h7D2F: out_word = 8'h00;
		16'h7D30: out_word = 8'hC9;
		16'h7D31: out_word = 8'hCD;
		16'h7D32: out_word = 8'h21;
		16'h7D33: out_word = 8'h3D;
		16'h7D34: out_word = 8'hE5;
		16'h7D35: out_word = 8'hC3;
		16'h7D36: out_word = 8'hF0;
		16'h7D37: out_word = 8'h3B;
		16'h7D38: out_word = 8'hAF;
		16'h7D39: out_word = 8'h00;
		16'h7D3A: out_word = 8'h00;
		16'h7D3B: out_word = 8'hDB;
		16'h7D3C: out_word = 8'hF7;
		16'h7D3D: out_word = 8'hFE;
		16'h7D3E: out_word = 8'h1E;
		16'h7D3F: out_word = 8'h28;
		16'h7D40: out_word = 8'h03;
		16'h7D41: out_word = 8'hFE;
		16'h7D42: out_word = 8'h1F;
		16'h7D43: out_word = 8'hC0;
		16'h7D44: out_word = 8'hCF;
		16'h7D45: out_word = 8'h31;
		16'h7D46: out_word = 8'h3E;
		16'h7D47: out_word = 8'h01;
		16'h7D48: out_word = 8'h32;
		16'h7D49: out_word = 8'hEF;
		16'h7D4A: out_word = 8'h5C;
		16'h7D4B: out_word = 8'hC9;
		16'h7D4C: out_word = 8'hAF;
		16'h7D4D: out_word = 8'hD3;
		16'h7D4E: out_word = 8'hFF;
		16'h7D4F: out_word = 8'hDB;
		16'h7D50: out_word = 8'hF6;
		16'h7D51: out_word = 8'h21;
		16'h7D52: out_word = 8'h38;
		16'h7D53: out_word = 8'h3D;
		16'h7D54: out_word = 8'h11;
		16'h7D55: out_word = 8'h92;
		16'h7D56: out_word = 8'h5C;
		16'h7D57: out_word = 8'h01;
		16'h7D58: out_word = 8'h14;
		16'h7D59: out_word = 8'h00;
		16'h7D5A: out_word = 8'hED;
		16'h7D5B: out_word = 8'hB0;
		16'h7D5C: out_word = 8'h21;
		16'h7D5D: out_word = 8'h67;
		16'h7D5E: out_word = 8'h3D;
		16'h7D5F: out_word = 8'hE5;
		16'h7D60: out_word = 8'h21;
		16'h7D61: out_word = 8'h2F;
		16'h7D62: out_word = 8'h3D;
		16'h7D63: out_word = 8'hE5;
		16'h7D64: out_word = 8'hC3;
		16'h7D65: out_word = 8'h92;
		16'h7D66: out_word = 8'h5C;
		16'h7D67: out_word = 8'h21;
		16'h7D68: out_word = 8'h90;
		16'h7D69: out_word = 8'h2F;
		16'h7D6A: out_word = 8'hE5;
		16'h7D6B: out_word = 8'h21;
		16'h7D6C: out_word = 8'h2F;
		16'h7D6D: out_word = 8'h3D;
		16'h7D6E: out_word = 8'hE5;
		16'h7D6F: out_word = 8'h21;
		16'h7D70: out_word = 8'h55;
		16'h7D71: out_word = 8'h16;
		16'h7D72: out_word = 8'hE5;
		16'h7D73: out_word = 8'h21;
		16'h7D74: out_word = 8'hFF;
		16'h7D75: out_word = 8'h5B;
		16'h7D76: out_word = 8'hE5;
		16'h7D77: out_word = 8'h36;
		16'h7D78: out_word = 8'hC9;
		16'h7D79: out_word = 8'h21;
		16'h7D7A: out_word = 8'hB5;
		16'h7D7B: out_word = 8'h5C;
		16'h7D7C: out_word = 8'h01;
		16'h7D7D: out_word = 8'h70;
		16'h7D7E: out_word = 8'h00;
		16'h7D7F: out_word = 8'hC9;
		16'h7D80: out_word = 8'h3E;
		16'h7D81: out_word = 8'h0D;
		16'h7D82: out_word = 8'hC3;
		16'h7D83: out_word = 8'h05;
		16'h7D84: out_word = 8'h08;
		16'h7D85: out_word = 8'hFF;
		16'h7D86: out_word = 8'hFF;
		16'h7D87: out_word = 8'h00;
		16'h7D88: out_word = 8'h00;
		16'h7D89: out_word = 8'hC3;
		16'h7D8A: out_word = 8'h17;
		16'h7D8B: out_word = 8'h08;
		16'h7D8C: out_word = 8'hFF;
		16'h7D8D: out_word = 8'hFF;
		16'h7D8E: out_word = 8'hFF;
		16'h7D8F: out_word = 8'h00;
		16'h7D90: out_word = 8'h00;
		16'h7D91: out_word = 8'hFF;
		16'h7D92: out_word = 8'hFF;
		16'h7D93: out_word = 8'hFF;
		16'h7D94: out_word = 8'hE7;
		16'h7D95: out_word = 8'h10;
		16'h7D96: out_word = 8'h00;
		16'h7D97: out_word = 8'hC9;
		16'h7D98: out_word = 8'h3E;
		16'h7D99: out_word = 8'h08;
		16'h7D9A: out_word = 8'hD3;
		16'h7D9B: out_word = 8'h1F;
		16'h7D9C: out_word = 8'hE5;
		16'h7D9D: out_word = 8'hE7;
		16'h7D9E: out_word = 8'h54;
		16'h7D9F: out_word = 8'h1F;
		16'h7DA0: out_word = 8'h38;
		16'h7DA1: out_word = 8'h03;
		16'h7DA2: out_word = 8'hE7;
		16'h7DA3: out_word = 8'h7B;
		16'h7DA4: out_word = 8'h1B;
		16'h7DA5: out_word = 8'hE1;
		16'h7DA6: out_word = 8'hDB;
		16'h7DA7: out_word = 8'hFF;
		16'h7DA8: out_word = 8'hE6;
		16'h7DA9: out_word = 8'h80;
		16'h7DAA: out_word = 8'h28;
		16'h7DAB: out_word = 8'hF0;
		16'h7DAC: out_word = 8'hC9;
		16'h7DAD: out_word = 8'h3E;
		16'h7DAE: out_word = 8'h08;
		16'h7DAF: out_word = 8'hCD;
		16'h7DB0: out_word = 8'h9A;
		16'h7DB1: out_word = 8'h3D;
		16'h7DB2: out_word = 8'h11;
		16'h7DB3: out_word = 8'h00;
		16'h7DB4: out_word = 8'h00;
		16'h7DB5: out_word = 8'hDB;
		16'h7DB6: out_word = 8'h1F;
		16'h7DB7: out_word = 8'hE6;
		16'h7DB8: out_word = 8'h02;
		16'h7DB9: out_word = 8'h47;
		16'h7DBA: out_word = 8'hDB;
		16'h7DBB: out_word = 8'h1F;
		16'h7DBC: out_word = 8'hE6;
		16'h7DBD: out_word = 8'h02;
		16'h7DBE: out_word = 8'hB8;
		16'h7DBF: out_word = 8'hC0;
		16'h7DC0: out_word = 8'h13;
		16'h7DC1: out_word = 8'h7B;
		16'h7DC2: out_word = 8'hB2;
		16'h7DC3: out_word = 8'h20;
		16'h7DC4: out_word = 8'hF5;
		16'h7DC5: out_word = 8'hC3;
		16'h7DC6: out_word = 8'hE7;
		16'h7DC7: out_word = 8'h3E;
		16'h7DC8: out_word = 8'h3A;
		16'h7DC9: out_word = 8'h19;
		16'h7DCA: out_word = 8'h5D;
		16'h7DCB: out_word = 8'hC3;
		16'h7DCC: out_word = 8'h12;
		16'h7DCD: out_word = 8'h39;
		16'h7DCE: out_word = 8'h21;
		16'h7DCF: out_word = 8'h16;
		16'h7DD0: out_word = 8'h5D;
		16'h7DD1: out_word = 8'h4F;
		16'h7DD2: out_word = 8'h3E;
		16'h7DD3: out_word = 8'h3C;
		16'h7DD4: out_word = 8'hB1;
		16'h7DD5: out_word = 8'hD3;
		16'h7DD6: out_word = 8'hFF;
		16'h7DD7: out_word = 8'h77;
		16'h7DD8: out_word = 8'hCD;
		16'h7DD9: out_word = 8'h08;
		16'h7DDA: out_word = 8'h3E;
		16'h7DDB: out_word = 8'hE6;
		16'h7DDC: out_word = 8'h80;
		16'h7DDD: out_word = 8'h28;
		16'h7DDE: out_word = 8'h1B;
		16'h7DDF: out_word = 8'hCD;
		16'h7DE0: out_word = 8'hAD;
		16'h7DE1: out_word = 8'h3D;
		16'h7DE2: out_word = 8'hCD;
		16'h7DE3: out_word = 8'h16;
		16'h7DE4: out_word = 8'h3E;
		16'h7DE5: out_word = 8'hCD;
		16'h7DE6: out_word = 8'h11;
		16'h7DE7: out_word = 8'h3E;
		16'h7DE8: out_word = 8'hFE;
		16'h7DE9: out_word = 8'hFF;
		16'h7DEA: out_word = 8'h20;
		16'h7DEB: out_word = 8'h0E;
		16'h7DEC: out_word = 8'hE5;
		16'h7DED: out_word = 8'hCD;
		16'h7DEE: out_word = 8'hCA;
		16'h7DEF: out_word = 8'h1F;
		16'h7DF0: out_word = 8'hE1;
		16'h7DF1: out_word = 8'hFE;
		16'h7DF2: out_word = 8'h50;
		16'h7DF3: out_word = 8'h3E;
		16'h7DF4: out_word = 8'h00;
		16'h7DF5: out_word = 8'h20;
		16'h7DF6: out_word = 8'h02;
		16'h7DF7: out_word = 8'h3E;
		16'h7DF8: out_word = 8'h80;
		16'h7DF9: out_word = 8'h77;
		16'h7DFA: out_word = 8'hCD;
		16'h7DFB: out_word = 8'h36;
		16'h7DFC: out_word = 8'h1E;
		16'h7DFD: out_word = 8'h3E;
		16'h7DFE: out_word = 8'h50;
		16'h7DFF: out_word = 8'h0E;
		16'h7E00: out_word = 8'hFF;
		16'h7E01: out_word = 8'h0D;
		16'h7E02: out_word = 8'h20;
		16'h7E03: out_word = 8'hFD;
		16'h7E04: out_word = 8'h3D;
		16'h7E05: out_word = 8'h20;
		16'h7E06: out_word = 8'hF8;
		16'h7E07: out_word = 8'hC9;
		16'h7E08: out_word = 8'h11;
		16'h7E09: out_word = 8'hFA;
		16'h7E0A: out_word = 8'h5C;
		16'h7E0B: out_word = 8'h2A;
		16'h7E0C: out_word = 8'hF6;
		16'h7E0D: out_word = 8'h5C;
		16'h7E0E: out_word = 8'h19;
		16'h7E0F: out_word = 8'h7E;
		16'h7E10: out_word = 8'hC9;
		16'h7E11: out_word = 8'h11;
		16'h7E12: out_word = 8'hC8;
		16'h7E13: out_word = 8'h5C;
		16'h7E14: out_word = 8'h18;
		16'h7E15: out_word = 8'hF5;
		16'h7E16: out_word = 8'hCD;
		16'h7E17: out_word = 8'h08;
		16'h7E18: out_word = 8'h3E;
		16'h7E19: out_word = 8'h06;
		16'h7E1A: out_word = 8'h08;
		16'h7E1B: out_word = 8'h0E;
		16'h7E1C: out_word = 8'h04;
		16'h7E1D: out_word = 8'h70;
		16'h7E1E: out_word = 8'h3E;
		16'h7E1F: out_word = 8'h08;
		16'h7E20: out_word = 8'hCD;
		16'h7E21: out_word = 8'h9A;
		16'h7E22: out_word = 8'h3D;
		16'h7E23: out_word = 8'hC9;
		16'h7E24: out_word = 8'h10;
		16'h7E25: out_word = 8'h06;
		16'h7E26: out_word = 8'h0B;
		16'h7E27: out_word = 8'hCD;
		16'h7E28: out_word = 8'h44;
		16'h7E29: out_word = 8'h3E;
		16'h7E2A: out_word = 8'h46;
		16'h7E2B: out_word = 8'h3E;
		16'h7E2C: out_word = 8'h01;
		16'h7E2D: out_word = 8'hCD;
		16'h7E2E: out_word = 8'h44;
		16'h7E2F: out_word = 8'h3E;
		16'h7E30: out_word = 8'hDB;
		16'h7E31: out_word = 8'h1F;
		16'h7E32: out_word = 8'hE6;
		16'h7E33: out_word = 8'h04;
		16'h7E34: out_word = 8'h20;
		16'h7E35: out_word = 8'h09;
		16'h7E36: out_word = 8'hAF;
		16'h7E37: out_word = 8'hCD;
		16'h7E38: out_word = 8'h44;
		16'h7E39: out_word = 8'h3E;
		16'h7E3A: out_word = 8'hDB;
		16'h7E3B: out_word = 8'h1F;
		16'h7E3C: out_word = 8'hE6;
		16'h7E3D: out_word = 8'h04;
		16'h7E3E: out_word = 8'hC0;
		16'h7E3F: out_word = 8'h04;
		16'h7E40: out_word = 8'h0D;
		16'h7E41: out_word = 8'hC8;
		16'h7E42: out_word = 8'h18;
		16'h7E43: out_word = 8'hD9;
		16'h7E44: out_word = 8'hD3;
		16'h7E45: out_word = 8'h7F;
		16'h7E46: out_word = 8'h78;
		16'h7E47: out_word = 8'hF6;
		16'h7E48: out_word = 8'h18;
		16'h7E49: out_word = 8'hC3;
		16'h7E4A: out_word = 8'h00;
		16'h7E4B: out_word = 8'h08;
		16'h7E4C: out_word = 8'hD3;
		16'h7E4D: out_word = 8'h7F;
		16'h7E4E: out_word = 8'hC3;
		16'h7E4F: out_word = 8'h80;
		16'h7E50: out_word = 8'h37;
		16'h7E51: out_word = 8'h3F;
		16'h7E52: out_word = 8'hB8;
		16'h7E53: out_word = 8'hC1;
		16'h7E54: out_word = 8'hF5;
		16'h7E55: out_word = 8'h78;
		16'h7E56: out_word = 8'hF6;
		16'h7E57: out_word = 8'h18;
		16'h7E58: out_word = 8'hCD;
		16'h7E59: out_word = 8'h00;
		16'h7E5A: out_word = 8'h08;
		16'h7E5B: out_word = 8'hF1;
		16'h7E5C: out_word = 8'hC8;
		16'h7E5D: out_word = 8'hC5;
		16'h7E5E: out_word = 8'hCD;
		16'h7E5F: out_word = 8'hFD;
		16'h7E60: out_word = 8'h3D;
		16'h7E61: out_word = 8'hC1;
		16'h7E62: out_word = 8'hC9;
		16'h7E63: out_word = 8'h4F;
		16'h7E64: out_word = 8'hCD;
		16'h7E65: out_word = 8'hEB;
		16'h7E66: out_word = 8'h1F;
		16'h7E67: out_word = 8'hCD;
		16'h7E68: out_word = 8'h11;
		16'h7E69: out_word = 8'h3E;
		16'h7E6A: out_word = 8'hE6;
		16'h7E6B: out_word = 8'h02;
		16'h7E6C: out_word = 8'hC4;
		16'h7E6D: out_word = 8'hAA;
		16'h7E6E: out_word = 8'h3E;
		16'h7E6F: out_word = 8'hC5;
		16'h7E70: out_word = 8'hCB;
		16'h7E71: out_word = 8'h7E;
		16'h7E72: out_word = 8'h28;
		16'h7E73: out_word = 8'h0F;
		16'h7E74: out_word = 8'hCB;
		16'h7E75: out_word = 8'h46;
		16'h7E76: out_word = 8'h20;
		16'h7E77: out_word = 8'h0B;
		16'h7E78: out_word = 8'hDB;
		16'h7E79: out_word = 8'h3F;
		16'h7E7A: out_word = 8'hB9;
		16'h7E7B: out_word = 8'h28;
		16'h7E7C: out_word = 8'h05;
		16'h7E7D: out_word = 8'h07;
		16'h7E7E: out_word = 8'hD3;
		16'h7E7F: out_word = 8'h3F;
		16'h7E80: out_word = 8'h79;
		16'h7E81: out_word = 8'h07;
		16'h7E82: out_word = 8'h4F;
		16'h7E83: out_word = 8'hCD;
		16'h7E84: out_word = 8'h08;
		16'h7E85: out_word = 8'h3E;
		16'h7E86: out_word = 8'h47;
		16'h7E87: out_word = 8'hDB;
		16'h7E88: out_word = 8'h3F;
		16'h7E89: out_word = 8'hB9;
		16'h7E8A: out_word = 8'hC5;
		16'h7E8B: out_word = 8'hC4;
		16'h7E8C: out_word = 8'h30;
		16'h7E8D: out_word = 8'h3D;
		16'h7E8E: out_word = 8'hC1;
		16'h7E8F: out_word = 8'h79;
		16'h7E90: out_word = 8'hCD;
		16'h7E91: out_word = 8'h4C;
		16'h7E92: out_word = 8'h3E;
		16'h7E93: out_word = 8'hC1;
		16'h7E94: out_word = 8'h79;
		16'h7E95: out_word = 8'hD3;
		16'h7E96: out_word = 8'h3F;
		16'h7E97: out_word = 8'h3A;
		16'h7E98: out_word = 8'hCD;
		16'h7E99: out_word = 8'h5C;
		16'h7E9A: out_word = 8'hB7;
		16'h7E9B: out_word = 8'hC8;
		16'h7E9C: out_word = 8'hAF;
		16'h7E9D: out_word = 8'h32;
		16'h7E9E: out_word = 8'hCD;
		16'h7E9F: out_word = 8'h5C;
		16'h7EA0: out_word = 8'h06;
		16'h7EA1: out_word = 8'h03;
		16'h7EA2: out_word = 8'h3E;
		16'h7EA3: out_word = 8'hFF;
		16'h7EA4: out_word = 8'hCD;
		16'h7EA5: out_word = 8'hFF;
		16'h7EA6: out_word = 8'h3D;
		16'h7EA7: out_word = 8'h10;
		16'h7EA8: out_word = 8'hF9;
		16'h7EA9: out_word = 8'hC9;
		16'h7EAA: out_word = 8'h79;
		16'h7EAB: out_word = 8'hB7;
		16'h7EAC: out_word = 8'h1F;
		16'h7EAD: out_word = 8'h4F;
		16'h7EAE: out_word = 8'hD0;
		16'h7EAF: out_word = 8'hC3;
		16'h7EB0: out_word = 8'hF6;
		16'h7EB1: out_word = 8'h1F;
		16'h7EB2: out_word = 8'hCD;
		16'h7EB3: out_word = 8'hEB;
		16'h7EB4: out_word = 8'h1F;
		16'h7EB5: out_word = 8'hDB;
		16'h7EB6: out_word = 8'h1F;
		16'h7EB7: out_word = 8'hE6;
		16'h7EB8: out_word = 8'h80;
		16'h7EB9: out_word = 8'h32;
		16'h7EBA: out_word = 8'hCD;
		16'h7EBB: out_word = 8'h5C;
		16'h7EBC: out_word = 8'hDB;
		16'h7EBD: out_word = 8'h3F;
		16'h7EBE: out_word = 8'h67;
		16'h7EBF: out_word = 8'hCD;
		16'h7EC0: out_word = 8'hCD;
		16'h7EC1: out_word = 8'h37;
		16'h7EC2: out_word = 8'h0E;
		16'h7EC3: out_word = 8'h7F;
		16'h7EC4: out_word = 8'h16;
		16'h7EC5: out_word = 8'h01;
		16'h7EC6: out_word = 8'hF3;
		16'h7EC7: out_word = 8'h3E;
		16'h7EC8: out_word = 8'hC0;
		16'h7EC9: out_word = 8'hD3;
		16'h7ECA: out_word = 8'h1F;
		16'h7ECB: out_word = 8'hC5;
		16'h7ECC: out_word = 8'h06;
		16'h7ECD: out_word = 8'h03;
		16'h7ECE: out_word = 8'hDB;
		16'h7ECF: out_word = 8'hFF;
		16'h7ED0: out_word = 8'hE6;
		16'h7ED1: out_word = 8'hC0;
		16'h7ED2: out_word = 8'h20;
		16'h7ED3: out_word = 8'h1E;
		16'h7ED4: out_word = 8'h13;
		16'h7ED5: out_word = 8'h7B;
		16'h7ED6: out_word = 8'hB2;
		16'h7ED7: out_word = 8'h20;
		16'h7ED8: out_word = 8'hF5;
		16'h7ED9: out_word = 8'h10;
		16'h7EDA: out_word = 8'hF3;
		16'h7EDB: out_word = 8'hC1;
		16'h7EDC: out_word = 8'hFB;
		16'h7EDD: out_word = 8'h3E;
		16'h7EDE: out_word = 8'hD0;
		16'h7EDF: out_word = 8'hD3;
		16'h7EE0: out_word = 8'h1F;
		16'h7EE1: out_word = 8'h3A;
		16'h7EE2: out_word = 8'hD1;
		16'h7EE3: out_word = 8'h5C;
		16'h7EE4: out_word = 8'hFE;
		16'h7EE5: out_word = 8'hFF;
		16'h7EE6: out_word = 8'hC8;
		16'h7EE7: out_word = 8'hCD;
		16'h7EE8: out_word = 8'h2B;
		16'h7EE9: out_word = 8'h27;
		16'h7EEA: out_word = 8'h3E;
		16'h7EEB: out_word = 8'hFF;
		16'h7EEC: out_word = 8'h32;
		16'h7EED: out_word = 8'h17;
		16'h7EEE: out_word = 8'h5D;
		16'h7EEF: out_word = 8'hC3;
		16'h7EF0: out_word = 8'h1B;
		16'h7EF1: out_word = 8'h27;
		16'h7EF2: out_word = 8'hC1;
		16'h7EF3: out_word = 8'hED;
		16'h7EF4: out_word = 8'h60;
		16'h7EF5: out_word = 8'hDB;
		16'h7EF6: out_word = 8'hFF;
		16'h7EF7: out_word = 8'hE6;
		16'h7EF8: out_word = 8'hC0;
		16'h7EF9: out_word = 8'h28;
		16'h7EFA: out_word = 8'hFA;
		16'h7EFB: out_word = 8'hFB;
		16'h7EFC: out_word = 8'hF8;
		16'h7EFD: out_word = 8'hF3;
		16'h7EFE: out_word = 8'hDB;
		16'h7EFF: out_word = 8'h7F;
		16'h7F00: out_word = 8'h18;
		16'h7F01: out_word = 8'hF3;
		16'h7F02: out_word = 8'h32;
		16'h7F03: out_word = 8'hFF;
		16'h7F04: out_word = 8'h5C;
		16'h7F05: out_word = 8'hC9;
		16'h7F06: out_word = 8'h22;
		16'h7F07: out_word = 8'h00;
		16'h7F08: out_word = 8'h5D;
		16'h7F09: out_word = 8'hC9;
		16'h7F0A: out_word = 8'h3E;
		16'h7F0B: out_word = 8'hA0;
		16'h7F0C: out_word = 8'h18;
		16'h7F0D: out_word = 8'h02;
		16'h7F0E: out_word = 8'h3E;
		16'h7F0F: out_word = 8'h80;
		16'h7F10: out_word = 8'h32;
		16'h7F11: out_word = 8'hFE;
		16'h7F12: out_word = 8'h5C;
		16'h7F13: out_word = 8'h16;
		16'h7F14: out_word = 8'h0A;
		16'h7F15: out_word = 8'hD5;
		16'h7F16: out_word = 8'hF3;
		16'h7F17: out_word = 8'h3A;
		16'h7F18: out_word = 8'hFF;
		16'h7F19: out_word = 8'h5C;
		16'h7F1A: out_word = 8'h3C;
		16'h7F1B: out_word = 8'hD3;
		16'h7F1C: out_word = 8'h5F;
		16'h7F1D: out_word = 8'h2A;
		16'h7F1E: out_word = 8'h00;
		16'h7F1F: out_word = 8'h5D;
		16'h7F20: out_word = 8'h0E;
		16'h7F21: out_word = 8'h7F;
		16'h7F22: out_word = 8'h3A;
		16'h7F23: out_word = 8'hFE;
		16'h7F24: out_word = 8'h5C;
		16'h7F25: out_word = 8'hD3;
		16'h7F26: out_word = 8'h1F;
		16'h7F27: out_word = 8'hFE;
		16'h7F28: out_word = 8'hA0;
		16'h7F29: out_word = 8'hF5;
		16'h7F2A: out_word = 8'hCC;
		16'h7F2B: out_word = 8'hBA;
		16'h7F2C: out_word = 8'h3F;
		16'h7F2D: out_word = 8'hF1;
		16'h7F2E: out_word = 8'hC4;
		16'h7F2F: out_word = 8'hD5;
		16'h7F30: out_word = 8'h3F;
		16'h7F31: out_word = 8'hD1;
		16'h7F32: out_word = 8'hFB;
		16'h7F33: out_word = 8'hDB;
		16'h7F34: out_word = 8'h1F;
		16'h7F35: out_word = 8'h47;
		16'h7F36: out_word = 8'hE6;
		16'h7F37: out_word = 8'h7F;
		16'h7F38: out_word = 8'hC8;
		16'h7F39: out_word = 8'h21;
		16'h7F3A: out_word = 8'hD8;
		16'h7F3B: out_word = 8'h29;
		16'h7F3C: out_word = 8'hE6;
		16'h7F3D: out_word = 8'h40;
		16'h7F3E: out_word = 8'h20;
		16'h7F3F: out_word = 8'h0B;
		16'h7F40: out_word = 8'h78;
		16'h7F41: out_word = 8'hE6;
		16'h7F42: out_word = 8'h04;
		16'h7F43: out_word = 8'h28;
		16'h7F44: out_word = 8'h5B;
		16'h7F45: out_word = 8'h15;
		16'h7F46: out_word = 8'h20;
		16'h7F47: out_word = 8'hCD;
		16'h7F48: out_word = 8'h21;
		16'h7F49: out_word = 8'hE2;
		16'h7F4A: out_word = 8'h29;
		16'h7F4B: out_word = 8'h3E;
		16'h7F4C: out_word = 8'hD0;
		16'h7F4D: out_word = 8'hD3;
		16'h7F4E: out_word = 8'h1F;
		16'h7F4F: out_word = 8'h78;
		16'h7F50: out_word = 8'hE6;
		16'h7F51: out_word = 8'h01;
		16'h7F52: out_word = 8'hC2;
		16'h7F53: out_word = 8'hE7;
		16'h7F54: out_word = 8'h3E;
		16'h7F55: out_word = 8'hDB;
		16'h7F56: out_word = 8'h3F;
		16'h7F57: out_word = 8'hB7;
		16'h7F58: out_word = 8'h20;
		16'h7F59: out_word = 8'h05;
		16'h7F5A: out_word = 8'hDB;
		16'h7F5B: out_word = 8'h5F;
		16'h7F5C: out_word = 8'hFE;
		16'h7F5D: out_word = 8'h0A;
		16'h7F5E: out_word = 8'hC8;
		16'h7F5F: out_word = 8'hE5;
		16'h7F60: out_word = 8'hCD;
		16'h7F61: out_word = 8'h97;
		16'h7F62: out_word = 8'h1D;
		16'h7F63: out_word = 8'hE1;
		16'h7F64: out_word = 8'hDF;
		16'h7F65: out_word = 8'h21;
		16'h7F66: out_word = 8'h13;
		16'h7F67: out_word = 8'h2A;
		16'h7F68: out_word = 8'hDF;
		16'h7F69: out_word = 8'hDB;
		16'h7F6A: out_word = 8'h3F;
		16'h7F6B: out_word = 8'hCD;
		16'h7F6C: out_word = 8'hA3;
		16'h7F6D: out_word = 8'h1D;
		16'h7F6E: out_word = 8'h21;
		16'h7F6F: out_word = 8'h18;
		16'h7F70: out_word = 8'h2A;
		16'h7F71: out_word = 8'hDF;
		16'h7F72: out_word = 8'hDB;
		16'h7F73: out_word = 8'h5F;
		16'h7F74: out_word = 8'hCD;
		16'h7F75: out_word = 8'hA3;
		16'h7F76: out_word = 8'h1D;
		16'h7F77: out_word = 8'h21;
		16'h7F78: out_word = 8'hFE;
		16'h7F79: out_word = 8'h29;
		16'h7F7A: out_word = 8'hDF;
		16'h7F7B: out_word = 8'hCD;
		16'h7F7C: out_word = 8'h52;
		16'h7F7D: out_word = 8'h10;
		16'h7F7E: out_word = 8'hFE;
		16'h7F7F: out_word = 8'h49;
		16'h7F80: out_word = 8'hC8;
		16'h7F81: out_word = 8'hFE;
		16'h7F82: out_word = 8'h52;
		16'h7F83: out_word = 8'h28;
		16'h7F84: out_word = 8'h0F;
		16'h7F85: out_word = 8'hFE;
		16'h7F86: out_word = 8'h41;
		16'h7F87: out_word = 8'h20;
		16'h7F88: out_word = 8'hF2;
		16'h7F89: out_word = 8'hCD;
		16'h7F8A: out_word = 8'h2B;
		16'h7F8B: out_word = 8'h27;
		16'h7F8C: out_word = 8'h3E;
		16'h7F8D: out_word = 8'h07;
		16'h7F8E: out_word = 8'h32;
		16'h7F8F: out_word = 8'h0F;
		16'h7F90: out_word = 8'h5D;
		16'h7F91: out_word = 8'hC3;
		16'h7F92: out_word = 8'hD3;
		16'h7F93: out_word = 8'h01;
		16'h7F94: out_word = 8'h3A;
		16'h7F95: out_word = 8'hF5;
		16'h7F96: out_word = 8'h5C;
		16'h7F97: out_word = 8'hCD;
		16'h7F98: out_word = 8'h63;
		16'h7F99: out_word = 8'h3E;
		16'h7F9A: out_word = 8'hCD;
		16'h7F9B: out_word = 8'hA0;
		16'h7F9C: out_word = 8'h3E;
		16'h7F9D: out_word = 8'hC3;
		16'h7F9E: out_word = 8'h13;
		16'h7F9F: out_word = 8'h3F;
		16'h7FA0: out_word = 8'h15;
		16'h7FA1: out_word = 8'hCA;
		16'h7FA2: out_word = 8'h48;
		16'h7FA3: out_word = 8'h3F;
		16'h7FA4: out_word = 8'hD5;
		16'h7FA5: out_word = 8'hCD;
		16'h7FA6: out_word = 8'h08;
		16'h7FA7: out_word = 8'h3E;
		16'h7FA8: out_word = 8'hE6;
		16'h7FA9: out_word = 8'h02;
		16'h7FAA: out_word = 8'h20;
		16'h7FAB: out_word = 8'h01;
		16'h7FAC: out_word = 8'h34;
		16'h7FAD: out_word = 8'hCD;
		16'h7FAE: out_word = 8'h98;
		16'h7FAF: out_word = 8'h3D;
		16'h7FB0: out_word = 8'h3A;
		16'h7FB1: out_word = 8'hF5;
		16'h7FB2: out_word = 8'h5C;
		16'h7FB3: out_word = 8'hCD;
		16'h7FB4: out_word = 8'h63;
		16'h7FB5: out_word = 8'h3E;
		16'h7FB6: out_word = 8'hD1;
		16'h7FB7: out_word = 8'hC3;
		16'h7FB8: out_word = 8'h15;
		16'h7FB9: out_word = 8'h3F;
		16'h7FBA: out_word = 8'h06;
		16'h7FBB: out_word = 8'h04;
		16'h7FBC: out_word = 8'hDB;
		16'h7FBD: out_word = 8'hFF;
		16'h7FBE: out_word = 8'hE6;
		16'h7FBF: out_word = 8'hC0;
		16'h7FC0: out_word = 8'h20;
		16'h7FC1: out_word = 8'h0F;
		16'h7FC2: out_word = 8'h13;
		16'h7FC3: out_word = 8'h7B;
		16'h7FC4: out_word = 8'hB2;
		16'h7FC5: out_word = 8'h20;
		16'h7FC6: out_word = 8'hF5;
		16'h7FC7: out_word = 8'h10;
		16'h7FC8: out_word = 8'hF3;
		16'h7FC9: out_word = 8'hC9;
		16'h7FCA: out_word = 8'hDB;
		16'h7FCB: out_word = 8'hFF;
		16'h7FCC: out_word = 8'hE6;
		16'h7FCD: out_word = 8'hC0;
		16'h7FCE: out_word = 8'h28;
		16'h7FCF: out_word = 8'hFA;
		16'h7FD0: out_word = 8'hF8;
		16'h7FD1: out_word = 8'hED;
		16'h7FD2: out_word = 8'hA3;
		16'h7FD3: out_word = 8'h18;
		16'h7FD4: out_word = 8'hF5;
		16'h7FD5: out_word = 8'h06;
		16'h7FD6: out_word = 8'h04;
		16'h7FD7: out_word = 8'hDB;
		16'h7FD8: out_word = 8'hFF;
		16'h7FD9: out_word = 8'hE6;
		16'h7FDA: out_word = 8'hC0;
		16'h7FDB: out_word = 8'h20;
		16'h7FDC: out_word = 8'h0F;
		16'h7FDD: out_word = 8'h13;
		16'h7FDE: out_word = 8'h7B;
		16'h7FDF: out_word = 8'hB2;
		16'h7FE0: out_word = 8'h20;
		16'h7FE1: out_word = 8'hF5;
		16'h7FE2: out_word = 8'h10;
		16'h7FE3: out_word = 8'hF3;
		16'h7FE4: out_word = 8'hC9;
		16'h7FE5: out_word = 8'hDB;
		16'h7FE6: out_word = 8'hFF;
		16'h7FE7: out_word = 8'hE6;
		16'h7FE8: out_word = 8'hC0;
		16'h7FE9: out_word = 8'h28;
		16'h7FEA: out_word = 8'hFA;
		16'h7FEB: out_word = 8'hF8;
		16'h7FEC: out_word = 8'hED;
		16'h7FED: out_word = 8'hA2;
		16'h7FEE: out_word = 8'h18;
		16'h7FEF: out_word = 8'hF5;
		16'h7FF0: out_word = 8'hED;
		16'h7FF1: out_word = 8'h79;
		16'h7FF2: out_word = 8'hC9;
		16'h7FF3: out_word = 8'hED;
		16'h7FF4: out_word = 8'h78;
		16'h7FF5: out_word = 8'hC9;
		16'h7FF6: out_word = 8'hFF;
		16'h7FF7: out_word = 8'hFF;
		16'h7FF8: out_word = 8'hFF;
		16'h7FF9: out_word = 8'hFF;
		16'h7FFA: out_word = 8'hFF;
		16'h7FFB: out_word = 8'hFF;
		16'h7FFC: out_word = 8'hFF;
		16'h7FFD: out_word = 8'hFF;
		16'h7FFE: out_word = 8'hFF;
		16'h7FFF: out_word = 8'hFF;
		16'h8000: out_word = 8'hF3;
		16'h8001: out_word = 8'h01;
		16'h8002: out_word = 8'h2B;
		16'h8003: out_word = 8'h69;
		16'h8004: out_word = 8'h0B;
		16'h8005: out_word = 8'h78;
		16'h8006: out_word = 8'hB1;
		16'h8007: out_word = 8'h20;
		16'h8008: out_word = 8'hFB;
		16'h8009: out_word = 8'hC3;
		16'h800A: out_word = 8'hC7;
		16'h800B: out_word = 8'h00;
		16'h800C: out_word = 8'h00;
		16'h800D: out_word = 8'h00;
		16'h800E: out_word = 8'h00;
		16'h800F: out_word = 8'h00;
		16'h8010: out_word = 8'hEF;
		16'h8011: out_word = 8'h10;
		16'h8012: out_word = 8'h00;
		16'h8013: out_word = 8'hC9;
		16'h8014: out_word = 8'h00;
		16'h8015: out_word = 8'h00;
		16'h8016: out_word = 8'h00;
		16'h8017: out_word = 8'h00;
		16'h8018: out_word = 8'hEF;
		16'h8019: out_word = 8'h18;
		16'h801A: out_word = 8'h00;
		16'h801B: out_word = 8'hC9;
		16'h801C: out_word = 8'h00;
		16'h801D: out_word = 8'h00;
		16'h801E: out_word = 8'h00;
		16'h801F: out_word = 8'h00;
		16'h8020: out_word = 8'hEF;
		16'h8021: out_word = 8'h20;
		16'h8022: out_word = 8'h00;
		16'h8023: out_word = 8'hC9;
		16'h8024: out_word = 8'h00;
		16'h8025: out_word = 8'h00;
		16'h8026: out_word = 8'h00;
		16'h8027: out_word = 8'h00;
		16'h8028: out_word = 8'hE3;
		16'h8029: out_word = 8'hF5;
		16'h802A: out_word = 8'h7E;
		16'h802B: out_word = 8'h23;
		16'h802C: out_word = 8'h23;
		16'h802D: out_word = 8'h22;
		16'h802E: out_word = 8'h5A;
		16'h802F: out_word = 8'h5B;
		16'h8030: out_word = 8'h2B;
		16'h8031: out_word = 8'h66;
		16'h8032: out_word = 8'h6F;
		16'h8033: out_word = 8'hF1;
		16'h8034: out_word = 8'hC3;
		16'h8035: out_word = 8'h5C;
		16'h8036: out_word = 8'h00;
		16'h8037: out_word = 8'h00;
		16'h8038: out_word = 8'hE5;
		16'h8039: out_word = 8'h21;
		16'h803A: out_word = 8'h48;
		16'h803B: out_word = 8'h00;
		16'h803C: out_word = 8'hE5;
		16'h803D: out_word = 8'h21;
		16'h803E: out_word = 8'h00;
		16'h803F: out_word = 8'h5B;
		16'h8040: out_word = 8'hE5;
		16'h8041: out_word = 8'h21;
		16'h8042: out_word = 8'h38;
		16'h8043: out_word = 8'h00;
		16'h8044: out_word = 8'hE5;
		16'h8045: out_word = 8'hC3;
		16'h8046: out_word = 8'h00;
		16'h8047: out_word = 8'h5B;
		16'h8048: out_word = 8'hE1;
		16'h8049: out_word = 8'hC9;
		16'h804A: out_word = 8'h01;
		16'h804B: out_word = 8'hFD;
		16'h804C: out_word = 8'h7F;
		16'h804D: out_word = 8'hAF;
		16'h804E: out_word = 8'hF3;
		16'h804F: out_word = 8'hED;
		16'h8050: out_word = 8'h79;
		16'h8051: out_word = 8'h32;
		16'h8052: out_word = 8'h5C;
		16'h8053: out_word = 8'h5B;
		16'h8054: out_word = 8'hFB;
		16'h8055: out_word = 8'h3D;
		16'h8056: out_word = 8'hFD;
		16'h8057: out_word = 8'h77;
		16'h8058: out_word = 8'h00;
		16'h8059: out_word = 8'hC3;
		16'h805A: out_word = 8'h21;
		16'h805B: out_word = 8'h03;
		16'h805C: out_word = 8'h22;
		16'h805D: out_word = 8'h58;
		16'h805E: out_word = 8'h5B;
		16'h805F: out_word = 8'h21;
		16'h8060: out_word = 8'h14;
		16'h8061: out_word = 8'h5B;
		16'h8062: out_word = 8'hE3;
		16'h8063: out_word = 8'hE5;
		16'h8064: out_word = 8'h2A;
		16'h8065: out_word = 8'h58;
		16'h8066: out_word = 8'h5B;
		16'h8067: out_word = 8'hE3;
		16'h8068: out_word = 8'hC3;
		16'h8069: out_word = 8'h00;
		16'h806A: out_word = 8'h5B;
		16'h806B: out_word = 8'hF5;
		16'h806C: out_word = 8'hC5;
		16'h806D: out_word = 8'h01;
		16'h806E: out_word = 8'hFD;
		16'h806F: out_word = 8'h7F;
		16'h8070: out_word = 8'h3A;
		16'h8071: out_word = 8'h5C;
		16'h8072: out_word = 8'h5B;
		16'h8073: out_word = 8'hEE;
		16'h8074: out_word = 8'h10;
		16'h8075: out_word = 8'hF3;
		16'h8076: out_word = 8'h32;
		16'h8077: out_word = 8'h5C;
		16'h8078: out_word = 8'h5B;
		16'h8079: out_word = 8'hED;
		16'h807A: out_word = 8'h79;
		16'h807B: out_word = 8'hFB;
		16'h807C: out_word = 8'hC1;
		16'h807D: out_word = 8'hF1;
		16'h807E: out_word = 8'hC9;
		16'h807F: out_word = 8'hCD;
		16'h8080: out_word = 8'h00;
		16'h8081: out_word = 8'h5B;
		16'h8082: out_word = 8'hE5;
		16'h8083: out_word = 8'h2A;
		16'h8084: out_word = 8'h5A;
		16'h8085: out_word = 8'h5B;
		16'h8086: out_word = 8'hE3;
		16'h8087: out_word = 8'hC9;
		16'h8088: out_word = 8'hF3;
		16'h8089: out_word = 8'h3A;
		16'h808A: out_word = 8'h5C;
		16'h808B: out_word = 8'h5B;
		16'h808C: out_word = 8'hE6;
		16'h808D: out_word = 8'hEF;
		16'h808E: out_word = 8'h32;
		16'h808F: out_word = 8'h5C;
		16'h8090: out_word = 8'h5B;
		16'h8091: out_word = 8'h01;
		16'h8092: out_word = 8'hFD;
		16'h8093: out_word = 8'h7F;
		16'h8094: out_word = 8'hED;
		16'h8095: out_word = 8'h79;
		16'h8096: out_word = 8'hFB;
		16'h8097: out_word = 8'hC3;
		16'h8098: out_word = 8'hC3;
		16'h8099: out_word = 8'h00;
		16'h809A: out_word = 8'h21;
		16'h809B: out_word = 8'hD8;
		16'h809C: out_word = 8'h06;
		16'h809D: out_word = 8'h18;
		16'h809E: out_word = 8'h03;
		16'h809F: out_word = 8'h21;
		16'h80A0: out_word = 8'hCA;
		16'h80A1: out_word = 8'h07;
		16'h80A2: out_word = 8'h08;
		16'h80A3: out_word = 8'h01;
		16'h80A4: out_word = 8'hFD;
		16'h80A5: out_word = 8'h7F;
		16'h80A6: out_word = 8'h3A;
		16'h80A7: out_word = 8'h5C;
		16'h80A8: out_word = 8'h5B;
		16'h80A9: out_word = 8'hF5;
		16'h80AA: out_word = 8'hE6;
		16'h80AB: out_word = 8'hEF;
		16'h80AC: out_word = 8'hF3;
		16'h80AD: out_word = 8'h32;
		16'h80AE: out_word = 8'h5C;
		16'h80AF: out_word = 8'h5B;
		16'h80B0: out_word = 8'hED;
		16'h80B1: out_word = 8'h79;
		16'h80B2: out_word = 8'hC3;
		16'h80B3: out_word = 8'hE6;
		16'h80B4: out_word = 8'h05;
		16'h80B5: out_word = 8'h08;
		16'h80B6: out_word = 8'hF1;
		16'h80B7: out_word = 8'h01;
		16'h80B8: out_word = 8'hFD;
		16'h80B9: out_word = 8'h7F;
		16'h80BA: out_word = 8'hF3;
		16'h80BB: out_word = 8'h32;
		16'h80BC: out_word = 8'h5C;
		16'h80BD: out_word = 8'h5B;
		16'h80BE: out_word = 8'hED;
		16'h80BF: out_word = 8'h79;
		16'h80C0: out_word = 8'hFB;
		16'h80C1: out_word = 8'h08;
		16'h80C2: out_word = 8'hC9;
		16'h80C3: out_word = 8'h2A;
		16'h80C4: out_word = 8'h8B;
		16'h80C5: out_word = 8'h5B;
		16'h80C6: out_word = 8'hE9;
		16'h80C7: out_word = 8'h06;
		16'h80C8: out_word = 8'h08;
		16'h80C9: out_word = 8'h78;
		16'h80CA: out_word = 8'hD9;
		16'h80CB: out_word = 8'h3D;
		16'h80CC: out_word = 8'h01;
		16'h80CD: out_word = 8'hFD;
		16'h80CE: out_word = 8'h7F;
		16'h80CF: out_word = 8'hED;
		16'h80D0: out_word = 8'h79;
		16'h80D1: out_word = 8'h21;
		16'h80D2: out_word = 8'h00;
		16'h80D3: out_word = 8'hC0;
		16'h80D4: out_word = 8'h11;
		16'h80D5: out_word = 8'h01;
		16'h80D6: out_word = 8'hC0;
		16'h80D7: out_word = 8'h01;
		16'h80D8: out_word = 8'hFF;
		16'h80D9: out_word = 8'h3F;
		16'h80DA: out_word = 8'h3E;
		16'h80DB: out_word = 8'hFF;
		16'h80DC: out_word = 8'h77;
		16'h80DD: out_word = 8'hBE;
		16'h80DE: out_word = 8'h20;
		16'h80DF: out_word = 8'h51;
		16'h80E0: out_word = 8'hAF;
		16'h80E1: out_word = 8'h77;
		16'h80E2: out_word = 8'hBE;
		16'h80E3: out_word = 8'h20;
		16'h80E4: out_word = 8'h4C;
		16'h80E5: out_word = 8'hED;
		16'h80E6: out_word = 8'hB0;
		16'h80E7: out_word = 8'hD9;
		16'h80E8: out_word = 8'h10;
		16'h80E9: out_word = 8'hDF;
		16'h80EA: out_word = 8'h32;
		16'h80EB: out_word = 8'h88;
		16'h80EC: out_word = 8'h5B;
		16'h80ED: out_word = 8'h0E;
		16'h80EE: out_word = 8'hFD;
		16'h80EF: out_word = 8'h16;
		16'h80F0: out_word = 8'hFF;
		16'h80F1: out_word = 8'h1E;
		16'h80F2: out_word = 8'hBF;
		16'h80F3: out_word = 8'h42;
		16'h80F4: out_word = 8'h3E;
		16'h80F5: out_word = 8'h0E;
		16'h80F6: out_word = 8'hED;
		16'h80F7: out_word = 8'h79;
		16'h80F8: out_word = 8'h43;
		16'h80F9: out_word = 8'h3E;
		16'h80FA: out_word = 8'hFF;
		16'h80FB: out_word = 8'hED;
		16'h80FC: out_word = 8'h79;
		16'h80FD: out_word = 8'h18;
		16'h80FE: out_word = 8'h38;
		16'h80FF: out_word = 8'h00;
		16'h8100: out_word = 8'hC3;
		16'h8101: out_word = 8'hAF;
		16'h8102: out_word = 8'h17;
		16'h8103: out_word = 8'hC3;
		16'h8104: out_word = 8'h38;
		16'h8105: out_word = 8'h18;
		16'h8106: out_word = 8'hC3;
		16'h8107: out_word = 8'hCF;
		16'h8108: out_word = 8'h1E;
		16'h8109: out_word = 8'hC3;
		16'h810A: out_word = 8'h04;
		16'h810B: out_word = 8'h1F;
		16'h810C: out_word = 8'hC3;
		16'h810D: out_word = 8'h4A;
		16'h810E: out_word = 8'h00;
		16'h810F: out_word = 8'hC3;
		16'h8110: out_word = 8'hA2;
		16'h8111: out_word = 8'h03;
		16'h8112: out_word = 8'hC3;
		16'h8113: out_word = 8'h2A;
		16'h8114: out_word = 8'h18;
		16'h8115: out_word = 8'hC3;
		16'h8116: out_word = 8'hA8;
		16'h8117: out_word = 8'h18;
		16'h8118: out_word = 8'hC3;
		16'h8119: out_word = 8'h2D;
		16'h811A: out_word = 8'h01;
		16'h811B: out_word = 8'hC3;
		16'h811C: out_word = 8'h05;
		16'h811D: out_word = 8'h0A;
		16'h811E: out_word = 8'hC3;
		16'h811F: out_word = 8'hA3;
		16'h8120: out_word = 8'h11;
		16'h8121: out_word = 8'hC3;
		16'h8122: out_word = 8'hD8;
		16'h8123: out_word = 8'h06;
		16'h8124: out_word = 8'hC3;
		16'h8125: out_word = 8'hCA;
		16'h8126: out_word = 8'h07;
		16'h8127: out_word = 8'hC3;
		16'h8128: out_word = 8'hA3;
		16'h8129: out_word = 8'h08;
		16'h812A: out_word = 8'hC3;
		16'h812B: out_word = 8'hF0;
		16'h812C: out_word = 8'h08;
		16'h812D: out_word = 8'hEF;
		16'h812E: out_word = 8'h01;
		16'h812F: out_word = 8'h3B;
		16'h8130: out_word = 8'hC9;
		16'h8131: out_word = 8'hD9;
		16'h8132: out_word = 8'h78;
		16'h8133: out_word = 8'hD3;
		16'h8134: out_word = 8'hFE;
		16'h8135: out_word = 8'h18;
		16'h8136: out_word = 8'hFE;
		16'h8137: out_word = 8'h42;
		16'h8138: out_word = 8'h3E;
		16'h8139: out_word = 8'h07;
		16'h813A: out_word = 8'hED;
		16'h813B: out_word = 8'h79;
		16'h813C: out_word = 8'h43;
		16'h813D: out_word = 8'h3E;
		16'h813E: out_word = 8'hFF;
		16'h813F: out_word = 8'hED;
		16'h8140: out_word = 8'h79;
		16'h8141: out_word = 8'h11;
		16'h8142: out_word = 8'h00;
		16'h8143: out_word = 8'h5B;
		16'h8144: out_word = 8'h21;
		16'h8145: out_word = 8'h6B;
		16'h8146: out_word = 8'h00;
		16'h8147: out_word = 8'h01;
		16'h8148: out_word = 8'h58;
		16'h8149: out_word = 8'h00;
		16'h814A: out_word = 8'hED;
		16'h814B: out_word = 8'hB0;
		16'h814C: out_word = 8'h3E;
		16'h814D: out_word = 8'hCF;
		16'h814E: out_word = 8'h32;
		16'h814F: out_word = 8'h5D;
		16'h8150: out_word = 8'h5B;
		16'h8151: out_word = 8'h31;
		16'h8152: out_word = 8'hFF;
		16'h8153: out_word = 8'h5B;
		16'h8154: out_word = 8'h3E;
		16'h8155: out_word = 8'h04;
		16'h8156: out_word = 8'hCD;
		16'h8157: out_word = 8'h64;
		16'h8158: out_word = 8'h1C;
		16'h8159: out_word = 8'hDD;
		16'h815A: out_word = 8'h21;
		16'h815B: out_word = 8'hEC;
		16'h815C: out_word = 8'hEB;
		16'h815D: out_word = 8'hDD;
		16'h815E: out_word = 8'h22;
		16'h815F: out_word = 8'h83;
		16'h8160: out_word = 8'h5B;
		16'h8161: out_word = 8'hDD;
		16'h8162: out_word = 8'h36;
		16'h8163: out_word = 8'h0A;
		16'h8164: out_word = 8'h00;
		16'h8165: out_word = 8'hDD;
		16'h8166: out_word = 8'h36;
		16'h8167: out_word = 8'h0B;
		16'h8168: out_word = 8'hC0;
		16'h8169: out_word = 8'hDD;
		16'h816A: out_word = 8'h36;
		16'h816B: out_word = 8'h0C;
		16'h816C: out_word = 8'h00;
		16'h816D: out_word = 8'h21;
		16'h816E: out_word = 8'hEC;
		16'h816F: out_word = 8'h2B;
		16'h8170: out_word = 8'h3E;
		16'h8171: out_word = 8'h01;
		16'h8172: out_word = 8'h22;
		16'h8173: out_word = 8'h85;
		16'h8174: out_word = 8'h5B;
		16'h8175: out_word = 8'h32;
		16'h8176: out_word = 8'h87;
		16'h8177: out_word = 8'h5B;
		16'h8178: out_word = 8'h3E;
		16'h8179: out_word = 8'h05;
		16'h817A: out_word = 8'hCD;
		16'h817B: out_word = 8'h64;
		16'h817C: out_word = 8'h1C;
		16'h817D: out_word = 8'h21;
		16'h817E: out_word = 8'hFF;
		16'h817F: out_word = 8'hFF;
		16'h8180: out_word = 8'h22;
		16'h8181: out_word = 8'hB4;
		16'h8182: out_word = 8'h5C;
		16'h8183: out_word = 8'h11;
		16'h8184: out_word = 8'hAF;
		16'h8185: out_word = 8'h3E;
		16'h8186: out_word = 8'h01;
		16'h8187: out_word = 8'hA8;
		16'h8188: out_word = 8'h00;
		16'h8189: out_word = 8'hEB;
		16'h818A: out_word = 8'hEF;
		16'h818B: out_word = 8'h61;
		16'h818C: out_word = 8'h16;
		16'h818D: out_word = 8'hEB;
		16'h818E: out_word = 8'h23;
		16'h818F: out_word = 8'h22;
		16'h8190: out_word = 8'h7B;
		16'h8191: out_word = 8'h5C;
		16'h8192: out_word = 8'h2B;
		16'h8193: out_word = 8'h01;
		16'h8194: out_word = 8'h40;
		16'h8195: out_word = 8'h00;
		16'h8196: out_word = 8'hED;
		16'h8197: out_word = 8'h43;
		16'h8198: out_word = 8'h38;
		16'h8199: out_word = 8'h5C;
		16'h819A: out_word = 8'h22;
		16'h819B: out_word = 8'hB2;
		16'h819C: out_word = 8'h5C;
		16'h819D: out_word = 8'h21;
		16'h819E: out_word = 8'h00;
		16'h819F: out_word = 8'h3C;
		16'h81A0: out_word = 8'h22;
		16'h81A1: out_word = 8'h36;
		16'h81A2: out_word = 8'h5C;
		16'h81A3: out_word = 8'h2A;
		16'h81A4: out_word = 8'hB2;
		16'h81A5: out_word = 8'h5C;
		16'h81A6: out_word = 8'h23;
		16'h81A7: out_word = 8'hF9;
		16'h81A8: out_word = 8'hED;
		16'h81A9: out_word = 8'h56;
		16'h81AA: out_word = 8'hFD;
		16'h81AB: out_word = 8'h21;
		16'h81AC: out_word = 8'h3A;
		16'h81AD: out_word = 8'h5C;
		16'h81AE: out_word = 8'hFD;
		16'h81AF: out_word = 8'hCB;
		16'h81B0: out_word = 8'h01;
		16'h81B1: out_word = 8'hE6;
		16'h81B2: out_word = 8'hFB;
		16'h81B3: out_word = 8'h21;
		16'h81B4: out_word = 8'h0B;
		16'h81B5: out_word = 8'h00;
		16'h81B6: out_word = 8'h22;
		16'h81B7: out_word = 8'h5F;
		16'h81B8: out_word = 8'h5B;
		16'h81B9: out_word = 8'hAF;
		16'h81BA: out_word = 8'h32;
		16'h81BB: out_word = 8'h61;
		16'h81BC: out_word = 8'h5B;
		16'h81BD: out_word = 8'h32;
		16'h81BE: out_word = 8'h63;
		16'h81BF: out_word = 8'h5B;
		16'h81C0: out_word = 8'h32;
		16'h81C1: out_word = 8'h65;
		16'h81C2: out_word = 8'h5B;
		16'h81C3: out_word = 8'h21;
		16'h81C4: out_word = 8'h00;
		16'h81C5: out_word = 8'hEC;
		16'h81C6: out_word = 8'h22;
		16'h81C7: out_word = 8'h24;
		16'h81C8: out_word = 8'hFF;
		16'h81C9: out_word = 8'h3E;
		16'h81CA: out_word = 8'h50;
		16'h81CB: out_word = 8'h32;
		16'h81CC: out_word = 8'h64;
		16'h81CD: out_word = 8'h5B;
		16'h81CE: out_word = 8'h21;
		16'h81CF: out_word = 8'h0A;
		16'h81D0: out_word = 8'h00;
		16'h81D1: out_word = 8'h22;
		16'h81D2: out_word = 8'h94;
		16'h81D3: out_word = 8'h5B;
		16'h81D4: out_word = 8'h22;
		16'h81D5: out_word = 8'h96;
		16'h81D6: out_word = 8'h5B;
		16'h81D7: out_word = 8'h21;
		16'h81D8: out_word = 8'hB6;
		16'h81D9: out_word = 8'h5C;
		16'h81DA: out_word = 8'h22;
		16'h81DB: out_word = 8'h4F;
		16'h81DC: out_word = 8'h5C;
		16'h81DD: out_word = 8'h11;
		16'h81DE: out_word = 8'h89;
		16'h81DF: out_word = 8'h05;
		16'h81E0: out_word = 8'h01;
		16'h81E1: out_word = 8'h15;
		16'h81E2: out_word = 8'h00;
		16'h81E3: out_word = 8'hEB;
		16'h81E4: out_word = 8'hED;
		16'h81E5: out_word = 8'hB0;
		16'h81E6: out_word = 8'hEB;
		16'h81E7: out_word = 8'h2B;
		16'h81E8: out_word = 8'h22;
		16'h81E9: out_word = 8'h57;
		16'h81EA: out_word = 8'h5C;
		16'h81EB: out_word = 8'h23;
		16'h81EC: out_word = 8'h22;
		16'h81ED: out_word = 8'h53;
		16'h81EE: out_word = 8'h5C;
		16'h81EF: out_word = 8'h22;
		16'h81F0: out_word = 8'h4B;
		16'h81F1: out_word = 8'h5C;
		16'h81F2: out_word = 8'h36;
		16'h81F3: out_word = 8'h80;
		16'h81F4: out_word = 8'h23;
		16'h81F5: out_word = 8'h22;
		16'h81F6: out_word = 8'h59;
		16'h81F7: out_word = 8'h5C;
		16'h81F8: out_word = 8'h36;
		16'h81F9: out_word = 8'h0D;
		16'h81FA: out_word = 8'h23;
		16'h81FB: out_word = 8'h36;
		16'h81FC: out_word = 8'h80;
		16'h81FD: out_word = 8'h23;
		16'h81FE: out_word = 8'h22;
		16'h81FF: out_word = 8'h61;
		16'h8200: out_word = 8'h5C;
		16'h8201: out_word = 8'h22;
		16'h8202: out_word = 8'h63;
		16'h8203: out_word = 8'h5C;
		16'h8204: out_word = 8'h22;
		16'h8205: out_word = 8'h65;
		16'h8206: out_word = 8'h5C;
		16'h8207: out_word = 8'h3E;
		16'h8208: out_word = 8'h38;
		16'h8209: out_word = 8'h32;
		16'h820A: out_word = 8'h8D;
		16'h820B: out_word = 8'h5C;
		16'h820C: out_word = 8'h32;
		16'h820D: out_word = 8'h8F;
		16'h820E: out_word = 8'h5C;
		16'h820F: out_word = 8'h32;
		16'h8210: out_word = 8'h48;
		16'h8211: out_word = 8'h5C;
		16'h8212: out_word = 8'hAF;
		16'h8213: out_word = 8'h32;
		16'h8214: out_word = 8'h13;
		16'h8215: out_word = 8'hEC;
		16'h8216: out_word = 8'h3E;
		16'h8217: out_word = 8'h07;
		16'h8218: out_word = 8'hD3;
		16'h8219: out_word = 8'hFE;
		16'h821A: out_word = 8'h21;
		16'h821B: out_word = 8'h23;
		16'h821C: out_word = 8'h05;
		16'h821D: out_word = 8'h22;
		16'h821E: out_word = 8'h09;
		16'h821F: out_word = 8'h5C;
		16'h8220: out_word = 8'hFD;
		16'h8221: out_word = 8'h35;
		16'h8222: out_word = 8'hC6;
		16'h8223: out_word = 8'hFD;
		16'h8224: out_word = 8'h35;
		16'h8225: out_word = 8'hCA;
		16'h8226: out_word = 8'h21;
		16'h8227: out_word = 8'h9E;
		16'h8228: out_word = 8'h05;
		16'h8229: out_word = 8'h11;
		16'h822A: out_word = 8'h10;
		16'h822B: out_word = 8'h5C;
		16'h822C: out_word = 8'h01;
		16'h822D: out_word = 8'h0E;
		16'h822E: out_word = 8'h00;
		16'h822F: out_word = 8'hED;
		16'h8230: out_word = 8'hB0;
		16'h8231: out_word = 8'hFD;
		16'h8232: out_word = 8'hCB;
		16'h8233: out_word = 8'h01;
		16'h8234: out_word = 8'h8E;
		16'h8235: out_word = 8'hFD;
		16'h8236: out_word = 8'h36;
		16'h8237: out_word = 8'h00;
		16'h8238: out_word = 8'hFF;
		16'h8239: out_word = 8'hFD;
		16'h823A: out_word = 8'h36;
		16'h823B: out_word = 8'h31;
		16'h823C: out_word = 8'h02;
		16'h823D: out_word = 8'hEF;
		16'h823E: out_word = 8'h6B;
		16'h823F: out_word = 8'h0D;
		16'h8240: out_word = 8'hEF;
		16'h8241: out_word = 8'h04;
		16'h8242: out_word = 8'h3C;
		16'h8243: out_word = 8'h11;
		16'h8244: out_word = 8'h61;
		16'h8245: out_word = 8'h05;
		16'h8246: out_word = 8'hCD;
		16'h8247: out_word = 8'h7D;
		16'h8248: out_word = 8'h05;
		16'h8249: out_word = 8'hFD;
		16'h824A: out_word = 8'h36;
		16'h824B: out_word = 8'h31;
		16'h824C: out_word = 8'h02;
		16'h824D: out_word = 8'hFD;
		16'h824E: out_word = 8'hCB;
		16'h824F: out_word = 8'h02;
		16'h8250: out_word = 8'hEE;
		16'h8251: out_word = 8'h21;
		16'h8252: out_word = 8'hFF;
		16'h8253: out_word = 8'h5B;
		16'h8254: out_word = 8'h22;
		16'h8255: out_word = 8'h81;
		16'h8256: out_word = 8'h5B;
		16'h8257: out_word = 8'hCD;
		16'h8258: out_word = 8'h45;
		16'h8259: out_word = 8'h1F;
		16'h825A: out_word = 8'h3E;
		16'h825B: out_word = 8'h38;
		16'h825C: out_word = 8'h32;
		16'h825D: out_word = 8'h11;
		16'h825E: out_word = 8'hEC;
		16'h825F: out_word = 8'h32;
		16'h8260: out_word = 8'h0F;
		16'h8261: out_word = 8'hEC;
		16'h8262: out_word = 8'hCD;
		16'h8263: out_word = 8'h84;
		16'h8264: out_word = 8'h25;
		16'h8265: out_word = 8'hCD;
		16'h8266: out_word = 8'h20;
		16'h8267: out_word = 8'h1F;
		16'h8268: out_word = 8'hC3;
		16'h8269: out_word = 8'h9F;
		16'h826A: out_word = 8'h25;
		16'h826B: out_word = 8'h21;
		16'h826C: out_word = 8'h66;
		16'h826D: out_word = 8'h5B;
		16'h826E: out_word = 8'hCB;
		16'h826F: out_word = 8'hC6;
		16'h8270: out_word = 8'hFD;
		16'h8271: out_word = 8'h36;
		16'h8272: out_word = 8'h00;
		16'h8273: out_word = 8'hFF;
		16'h8274: out_word = 8'hFD;
		16'h8275: out_word = 8'h36;
		16'h8276: out_word = 8'h31;
		16'h8277: out_word = 8'h02;
		16'h8278: out_word = 8'h21;
		16'h8279: out_word = 8'h1D;
		16'h827A: out_word = 8'h5B;
		16'h827B: out_word = 8'hE5;
		16'h827C: out_word = 8'hED;
		16'h827D: out_word = 8'h73;
		16'h827E: out_word = 8'h3D;
		16'h827F: out_word = 8'h5C;
		16'h8280: out_word = 8'h21;
		16'h8281: out_word = 8'hBA;
		16'h8282: out_word = 8'h02;
		16'h8283: out_word = 8'h22;
		16'h8284: out_word = 8'h8B;
		16'h8285: out_word = 8'h5B;
		16'h8286: out_word = 8'hCD;
		16'h8287: out_word = 8'h8E;
		16'h8288: out_word = 8'h22;
		16'h8289: out_word = 8'hCD;
		16'h828A: out_word = 8'hCB;
		16'h828B: out_word = 8'h22;
		16'h828C: out_word = 8'hCA;
		16'h828D: out_word = 8'hF8;
		16'h828E: out_word = 8'h21;
		16'h828F: out_word = 8'hFE;
		16'h8290: out_word = 8'h28;
		16'h8291: out_word = 8'hCA;
		16'h8292: out_word = 8'hF8;
		16'h8293: out_word = 8'h21;
		16'h8294: out_word = 8'hFE;
		16'h8295: out_word = 8'h2D;
		16'h8296: out_word = 8'hCA;
		16'h8297: out_word = 8'hF8;
		16'h8298: out_word = 8'h21;
		16'h8299: out_word = 8'hFE;
		16'h829A: out_word = 8'h2B;
		16'h829B: out_word = 8'hCA;
		16'h829C: out_word = 8'hF8;
		16'h829D: out_word = 8'h21;
		16'h829E: out_word = 8'hCD;
		16'h829F: out_word = 8'hE0;
		16'h82A0: out_word = 8'h22;
		16'h82A1: out_word = 8'hCA;
		16'h82A2: out_word = 8'hF8;
		16'h82A3: out_word = 8'h21;
		16'h82A4: out_word = 8'hCD;
		16'h82A5: out_word = 8'h45;
		16'h82A6: out_word = 8'h1F;
		16'h82A7: out_word = 8'h3A;
		16'h82A8: out_word = 8'h0E;
		16'h82A9: out_word = 8'hEC;
		16'h82AA: out_word = 8'hCD;
		16'h82AB: out_word = 8'h20;
		16'h82AC: out_word = 8'h1F;
		16'h82AD: out_word = 8'hFE;
		16'h82AE: out_word = 8'h04;
		16'h82AF: out_word = 8'hC2;
		16'h82B0: out_word = 8'hAF;
		16'h82B1: out_word = 8'h17;
		16'h82B2: out_word = 8'hCD;
		16'h82B3: out_word = 8'h97;
		16'h82B4: out_word = 8'h22;
		16'h82B5: out_word = 8'hCA;
		16'h82B6: out_word = 8'hAF;
		16'h82B7: out_word = 8'h17;
		16'h82B8: out_word = 8'hE1;
		16'h82B9: out_word = 8'hC9;
		16'h82BA: out_word = 8'hFD;
		16'h82BB: out_word = 8'hCB;
		16'h82BC: out_word = 8'h00;
		16'h82BD: out_word = 8'h7E;
		16'h82BE: out_word = 8'h20;
		16'h82BF: out_word = 8'h01;
		16'h82C0: out_word = 8'hC9;
		16'h82C1: out_word = 8'h2A;
		16'h82C2: out_word = 8'h59;
		16'h82C3: out_word = 8'h5C;
		16'h82C4: out_word = 8'h22;
		16'h82C5: out_word = 8'h5D;
		16'h82C6: out_word = 8'h5C;
		16'h82C7: out_word = 8'hEF;
		16'h82C8: out_word = 8'hFB;
		16'h82C9: out_word = 8'h19;
		16'h82CA: out_word = 8'h78;
		16'h82CB: out_word = 8'hB1;
		16'h82CC: out_word = 8'hC2;
		16'h82CD: out_word = 8'hF7;
		16'h82CE: out_word = 8'h03;
		16'h82CF: out_word = 8'hDF;
		16'h82D0: out_word = 8'hFE;
		16'h82D1: out_word = 8'h0D;
		16'h82D2: out_word = 8'hC8;
		16'h82D3: out_word = 8'hCD;
		16'h82D4: out_word = 8'hEF;
		16'h82D5: out_word = 8'h21;
		16'h82D6: out_word = 8'hFD;
		16'h82D7: out_word = 8'hCB;
		16'h82D8: out_word = 8'h02;
		16'h82D9: out_word = 8'h76;
		16'h82DA: out_word = 8'h20;
		16'h82DB: out_word = 8'h03;
		16'h82DC: out_word = 8'hEF;
		16'h82DD: out_word = 8'h6E;
		16'h82DE: out_word = 8'h0D;
		16'h82DF: out_word = 8'hFD;
		16'h82E0: out_word = 8'hCB;
		16'h82E1: out_word = 8'h02;
		16'h82E2: out_word = 8'hB6;
		16'h82E3: out_word = 8'hCD;
		16'h82E4: out_word = 8'h45;
		16'h82E5: out_word = 8'h1F;
		16'h82E6: out_word = 8'h21;
		16'h82E7: out_word = 8'h0D;
		16'h82E8: out_word = 8'hEC;
		16'h82E9: out_word = 8'hCB;
		16'h82EA: out_word = 8'h76;
		16'h82EB: out_word = 8'h20;
		16'h82EC: out_word = 8'h07;
		16'h82ED: out_word = 8'h23;
		16'h82EE: out_word = 8'h7E;
		16'h82EF: out_word = 8'hFE;
		16'h82F0: out_word = 8'h00;
		16'h82F1: out_word = 8'hCC;
		16'h82F2: out_word = 8'h81;
		16'h82F3: out_word = 8'h38;
		16'h82F4: out_word = 8'hCD;
		16'h82F5: out_word = 8'h20;
		16'h82F6: out_word = 8'h1F;
		16'h82F7: out_word = 8'h21;
		16'h82F8: out_word = 8'h3C;
		16'h82F9: out_word = 8'h5C;
		16'h82FA: out_word = 8'hCB;
		16'h82FB: out_word = 8'h9E;
		16'h82FC: out_word = 8'h3E;
		16'h82FD: out_word = 8'h19;
		16'h82FE: out_word = 8'hFD;
		16'h82FF: out_word = 8'h96;
		16'h8300: out_word = 8'h4F;
		16'h8301: out_word = 8'h32;
		16'h8302: out_word = 8'h8C;
		16'h8303: out_word = 8'h5C;
		16'h8304: out_word = 8'hFD;
		16'h8305: out_word = 8'hCB;
		16'h8306: out_word = 8'h01;
		16'h8307: out_word = 8'hFE;
		16'h8308: out_word = 8'hFD;
		16'h8309: out_word = 8'h36;
		16'h830A: out_word = 8'h0A;
		16'h830B: out_word = 8'h01;
		16'h830C: out_word = 8'h21;
		16'h830D: out_word = 8'h00;
		16'h830E: out_word = 8'h3E;
		16'h830F: out_word = 8'hE5;
		16'h8310: out_word = 8'h21;
		16'h8311: out_word = 8'h1D;
		16'h8312: out_word = 8'h5B;
		16'h8313: out_word = 8'hE5;
		16'h8314: out_word = 8'hED;
		16'h8315: out_word = 8'h73;
		16'h8316: out_word = 8'h3D;
		16'h8317: out_word = 8'h5C;
		16'h8318: out_word = 8'h21;
		16'h8319: out_word = 8'h21;
		16'h831A: out_word = 8'h03;
		16'h831B: out_word = 8'h22;
		16'h831C: out_word = 8'h8B;
		16'h831D: out_word = 8'h5B;
		16'h831E: out_word = 8'hC3;
		16'h831F: out_word = 8'h38;
		16'h8320: out_word = 8'h18;
		16'h8321: out_word = 8'hED;
		16'h8322: out_word = 8'h7B;
		16'h8323: out_word = 8'hB2;
		16'h8324: out_word = 8'h5C;
		16'h8325: out_word = 8'h33;
		16'h8326: out_word = 8'h21;
		16'h8327: out_word = 8'hFF;
		16'h8328: out_word = 8'h5B;
		16'h8329: out_word = 8'h22;
		16'h832A: out_word = 8'h81;
		16'h832B: out_word = 8'h5B;
		16'h832C: out_word = 8'h76;
		16'h832D: out_word = 8'hFD;
		16'h832E: out_word = 8'hCB;
		16'h832F: out_word = 8'h01;
		16'h8330: out_word = 8'hAE;
		16'h8331: out_word = 8'h21;
		16'h8332: out_word = 8'h66;
		16'h8333: out_word = 8'h5B;
		16'h8334: out_word = 8'hCB;
		16'h8335: out_word = 8'h56;
		16'h8336: out_word = 8'h28;
		16'h8337: out_word = 8'h12;
		16'h8338: out_word = 8'hCD;
		16'h8339: out_word = 8'h45;
		16'h833A: out_word = 8'h1F;
		16'h833B: out_word = 8'hDD;
		16'h833C: out_word = 8'h2A;
		16'h833D: out_word = 8'h83;
		16'h833E: out_word = 8'h5B;
		16'h833F: out_word = 8'h01;
		16'h8340: out_word = 8'h14;
		16'h8341: out_word = 8'h00;
		16'h8342: out_word = 8'hDD;
		16'h8343: out_word = 8'h09;
		16'h8344: out_word = 8'hCD;
		16'h8345: out_word = 8'h56;
		16'h8346: out_word = 8'h1D;
		16'h8347: out_word = 8'hCD;
		16'h8348: out_word = 8'h20;
		16'h8349: out_word = 8'h1F;
		16'h834A: out_word = 8'h3A;
		16'h834B: out_word = 8'h3A;
		16'h834C: out_word = 8'h5C;
		16'h834D: out_word = 8'h3C;
		16'h834E: out_word = 8'hF5;
		16'h834F: out_word = 8'h21;
		16'h8350: out_word = 8'h00;
		16'h8351: out_word = 8'h00;
		16'h8352: out_word = 8'hFD;
		16'h8353: out_word = 8'h74;
		16'h8354: out_word = 8'h37;
		16'h8355: out_word = 8'hFD;
		16'h8356: out_word = 8'h74;
		16'h8357: out_word = 8'h26;
		16'h8358: out_word = 8'h22;
		16'h8359: out_word = 8'h0B;
		16'h835A: out_word = 8'h5C;
		16'h835B: out_word = 8'h21;
		16'h835C: out_word = 8'h01;
		16'h835D: out_word = 8'h00;
		16'h835E: out_word = 8'h22;
		16'h835F: out_word = 8'h16;
		16'h8360: out_word = 8'h5C;
		16'h8361: out_word = 8'hEF;
		16'h8362: out_word = 8'hB0;
		16'h8363: out_word = 8'h16;
		16'h8364: out_word = 8'hFD;
		16'h8365: out_word = 8'hCB;
		16'h8366: out_word = 8'h37;
		16'h8367: out_word = 8'hAE;
		16'h8368: out_word = 8'hEF;
		16'h8369: out_word = 8'h6E;
		16'h836A: out_word = 8'h0D;
		16'h836B: out_word = 8'hFD;
		16'h836C: out_word = 8'hCB;
		16'h836D: out_word = 8'h02;
		16'h836E: out_word = 8'hEE;
		16'h836F: out_word = 8'hF1;
		16'h8370: out_word = 8'h47;
		16'h8371: out_word = 8'hFE;
		16'h8372: out_word = 8'h0A;
		16'h8373: out_word = 8'h38;
		16'h8374: out_word = 8'h0A;
		16'h8375: out_word = 8'hFE;
		16'h8376: out_word = 8'h1D;
		16'h8377: out_word = 8'h38;
		16'h8378: out_word = 8'h04;
		16'h8379: out_word = 8'hC6;
		16'h837A: out_word = 8'h14;
		16'h837B: out_word = 8'h18;
		16'h837C: out_word = 8'h02;
		16'h837D: out_word = 8'hC6;
		16'h837E: out_word = 8'h07;
		16'h837F: out_word = 8'hEF;
		16'h8380: out_word = 8'hEF;
		16'h8381: out_word = 8'h15;
		16'h8382: out_word = 8'h3E;
		16'h8383: out_word = 8'h20;
		16'h8384: out_word = 8'hD7;
		16'h8385: out_word = 8'h78;
		16'h8386: out_word = 8'hFE;
		16'h8387: out_word = 8'h1D;
		16'h8388: out_word = 8'h38;
		16'h8389: out_word = 8'h12;
		16'h838A: out_word = 8'hD6;
		16'h838B: out_word = 8'h1D;
		16'h838C: out_word = 8'h06;
		16'h838D: out_word = 8'h00;
		16'h838E: out_word = 8'h4F;
		16'h838F: out_word = 8'h21;
		16'h8390: out_word = 8'h6C;
		16'h8391: out_word = 8'h04;
		16'h8392: out_word = 8'h09;
		16'h8393: out_word = 8'h09;
		16'h8394: out_word = 8'h5E;
		16'h8395: out_word = 8'h23;
		16'h8396: out_word = 8'h56;
		16'h8397: out_word = 8'hCD;
		16'h8398: out_word = 8'h7D;
		16'h8399: out_word = 8'h05;
		16'h839A: out_word = 8'h18;
		16'h839B: out_word = 8'h06;
		16'h839C: out_word = 8'h11;
		16'h839D: out_word = 8'h91;
		16'h839E: out_word = 8'h13;
		16'h839F: out_word = 8'hEF;
		16'h83A0: out_word = 8'h0A;
		16'h83A1: out_word = 8'h0C;
		16'h83A2: out_word = 8'hAF;
		16'h83A3: out_word = 8'h11;
		16'h83A4: out_word = 8'h36;
		16'h83A5: out_word = 8'h15;
		16'h83A6: out_word = 8'hEF;
		16'h83A7: out_word = 8'h0A;
		16'h83A8: out_word = 8'h0C;
		16'h83A9: out_word = 8'hED;
		16'h83AA: out_word = 8'h4B;
		16'h83AB: out_word = 8'h45;
		16'h83AC: out_word = 8'h5C;
		16'h83AD: out_word = 8'hEF;
		16'h83AE: out_word = 8'h1B;
		16'h83AF: out_word = 8'h1A;
		16'h83B0: out_word = 8'h3E;
		16'h83B1: out_word = 8'h3A;
		16'h83B2: out_word = 8'hD7;
		16'h83B3: out_word = 8'hFD;
		16'h83B4: out_word = 8'h4E;
		16'h83B5: out_word = 8'h0D;
		16'h83B6: out_word = 8'h06;
		16'h83B7: out_word = 8'h00;
		16'h83B8: out_word = 8'hEF;
		16'h83B9: out_word = 8'h1B;
		16'h83BA: out_word = 8'h1A;
		16'h83BB: out_word = 8'hEF;
		16'h83BC: out_word = 8'h97;
		16'h83BD: out_word = 8'h10;
		16'h83BE: out_word = 8'h3A;
		16'h83BF: out_word = 8'h3A;
		16'h83C0: out_word = 8'h5C;
		16'h83C1: out_word = 8'h3C;
		16'h83C2: out_word = 8'h28;
		16'h83C3: out_word = 8'h1B;
		16'h83C4: out_word = 8'hFE;
		16'h83C5: out_word = 8'h09;
		16'h83C6: out_word = 8'h28;
		16'h83C7: out_word = 8'h04;
		16'h83C8: out_word = 8'hFE;
		16'h83C9: out_word = 8'h15;
		16'h83CA: out_word = 8'h20;
		16'h83CB: out_word = 8'h03;
		16'h83CC: out_word = 8'hFD;
		16'h83CD: out_word = 8'h34;
		16'h83CE: out_word = 8'h0D;
		16'h83CF: out_word = 8'h01;
		16'h83D0: out_word = 8'h03;
		16'h83D1: out_word = 8'h00;
		16'h83D2: out_word = 8'h11;
		16'h83D3: out_word = 8'h70;
		16'h83D4: out_word = 8'h5C;
		16'h83D5: out_word = 8'h21;
		16'h83D6: out_word = 8'h44;
		16'h83D7: out_word = 8'h5C;
		16'h83D8: out_word = 8'hCB;
		16'h83D9: out_word = 8'h7E;
		16'h83DA: out_word = 8'h28;
		16'h83DB: out_word = 8'h01;
		16'h83DC: out_word = 8'h09;
		16'h83DD: out_word = 8'hED;
		16'h83DE: out_word = 8'hB8;
		16'h83DF: out_word = 8'hFD;
		16'h83E0: out_word = 8'h36;
		16'h83E1: out_word = 8'h0A;
		16'h83E2: out_word = 8'hFF;
		16'h83E3: out_word = 8'hFD;
		16'h83E4: out_word = 8'hCB;
		16'h83E5: out_word = 8'h01;
		16'h83E6: out_word = 8'h9E;
		16'h83E7: out_word = 8'h21;
		16'h83E8: out_word = 8'h66;
		16'h83E9: out_word = 8'h5B;
		16'h83EA: out_word = 8'hCB;
		16'h83EB: out_word = 8'h86;
		16'h83EC: out_word = 8'hC3;
		16'h83ED: out_word = 8'hCB;
		16'h83EE: out_word = 8'h25;
		16'h83EF: out_word = 8'h3E;
		16'h83F0: out_word = 8'h10;
		16'h83F1: out_word = 8'h01;
		16'h83F2: out_word = 8'h00;
		16'h83F3: out_word = 8'h00;
		16'h83F4: out_word = 8'hC3;
		16'h83F5: out_word = 8'h4E;
		16'h83F6: out_word = 8'h03;
		16'h83F7: out_word = 8'hED;
		16'h83F8: out_word = 8'h43;
		16'h83F9: out_word = 8'h49;
		16'h83FA: out_word = 8'h5C;
		16'h83FB: out_word = 8'hCD;
		16'h83FC: out_word = 8'h45;
		16'h83FD: out_word = 8'h1F;
		16'h83FE: out_word = 8'h78;
		16'h83FF: out_word = 8'hB1;
		16'h8400: out_word = 8'h28;
		16'h8401: out_word = 8'h08;
		16'h8402: out_word = 8'hED;
		16'h8403: out_word = 8'h43;
		16'h8404: out_word = 8'h49;
		16'h8405: out_word = 8'h5C;
		16'h8406: out_word = 8'hED;
		16'h8407: out_word = 8'h43;
		16'h8408: out_word = 8'h08;
		16'h8409: out_word = 8'hEC;
		16'h840A: out_word = 8'hCD;
		16'h840B: out_word = 8'h20;
		16'h840C: out_word = 8'h1F;
		16'h840D: out_word = 8'h2A;
		16'h840E: out_word = 8'h5D;
		16'h840F: out_word = 8'h5C;
		16'h8410: out_word = 8'hEB;
		16'h8411: out_word = 8'h21;
		16'h8412: out_word = 8'hEF;
		16'h8413: out_word = 8'h03;
		16'h8414: out_word = 8'hE5;
		16'h8415: out_word = 8'h2A;
		16'h8416: out_word = 8'h61;
		16'h8417: out_word = 8'h5C;
		16'h8418: out_word = 8'h37;
		16'h8419: out_word = 8'hED;
		16'h841A: out_word = 8'h52;
		16'h841B: out_word = 8'hE5;
		16'h841C: out_word = 8'h60;
		16'h841D: out_word = 8'h69;
		16'h841E: out_word = 8'hEF;
		16'h841F: out_word = 8'h6E;
		16'h8420: out_word = 8'h19;
		16'h8421: out_word = 8'h20;
		16'h8422: out_word = 8'h06;
		16'h8423: out_word = 8'hEF;
		16'h8424: out_word = 8'hB8;
		16'h8425: out_word = 8'h19;
		16'h8426: out_word = 8'hEF;
		16'h8427: out_word = 8'hE8;
		16'h8428: out_word = 8'h19;
		16'h8429: out_word = 8'hC1;
		16'h842A: out_word = 8'h79;
		16'h842B: out_word = 8'h3D;
		16'h842C: out_word = 8'hB0;
		16'h842D: out_word = 8'h20;
		16'h842E: out_word = 8'h13;
		16'h842F: out_word = 8'hCD;
		16'h8430: out_word = 8'h45;
		16'h8431: out_word = 8'h1F;
		16'h8432: out_word = 8'hE5;
		16'h8433: out_word = 8'h2A;
		16'h8434: out_word = 8'h49;
		16'h8435: out_word = 8'h5C;
		16'h8436: out_word = 8'hCD;
		16'h8437: out_word = 8'h4A;
		16'h8438: out_word = 8'h33;
		16'h8439: out_word = 8'h22;
		16'h843A: out_word = 8'h49;
		16'h843B: out_word = 8'h5C;
		16'h843C: out_word = 8'hE1;
		16'h843D: out_word = 8'hCD;
		16'h843E: out_word = 8'h20;
		16'h843F: out_word = 8'h1F;
		16'h8440: out_word = 8'h18;
		16'h8441: out_word = 8'h28;
		16'h8442: out_word = 8'hC5;
		16'h8443: out_word = 8'h03;
		16'h8444: out_word = 8'h03;
		16'h8445: out_word = 8'h03;
		16'h8446: out_word = 8'h03;
		16'h8447: out_word = 8'h2B;
		16'h8448: out_word = 8'hED;
		16'h8449: out_word = 8'h5B;
		16'h844A: out_word = 8'h53;
		16'h844B: out_word = 8'h5C;
		16'h844C: out_word = 8'hD5;
		16'h844D: out_word = 8'hEF;
		16'h844E: out_word = 8'h55;
		16'h844F: out_word = 8'h16;
		16'h8450: out_word = 8'hE1;
		16'h8451: out_word = 8'h22;
		16'h8452: out_word = 8'h53;
		16'h8453: out_word = 8'h5C;
		16'h8454: out_word = 8'hC1;
		16'h8455: out_word = 8'hC5;
		16'h8456: out_word = 8'h13;
		16'h8457: out_word = 8'h2A;
		16'h8458: out_word = 8'h61;
		16'h8459: out_word = 8'h5C;
		16'h845A: out_word = 8'h2B;
		16'h845B: out_word = 8'h2B;
		16'h845C: out_word = 8'hED;
		16'h845D: out_word = 8'hB8;
		16'h845E: out_word = 8'h2A;
		16'h845F: out_word = 8'h49;
		16'h8460: out_word = 8'h5C;
		16'h8461: out_word = 8'hEB;
		16'h8462: out_word = 8'hC1;
		16'h8463: out_word = 8'h70;
		16'h8464: out_word = 8'h2B;
		16'h8465: out_word = 8'h71;
		16'h8466: out_word = 8'h2B;
		16'h8467: out_word = 8'h73;
		16'h8468: out_word = 8'h2B;
		16'h8469: out_word = 8'h72;
		16'h846A: out_word = 8'hF1;
		16'h846B: out_word = 8'hC9;
		16'h846C: out_word = 8'h8C;
		16'h846D: out_word = 8'h04;
		16'h846E: out_word = 8'h97;
		16'h846F: out_word = 8'h04;
		16'h8470: out_word = 8'hA6;
		16'h8471: out_word = 8'h04;
		16'h8472: out_word = 8'hB0;
		16'h8473: out_word = 8'h04;
		16'h8474: out_word = 8'hC1;
		16'h8475: out_word = 8'h04;
		16'h8476: out_word = 8'hD4;
		16'h8477: out_word = 8'h04;
		16'h8478: out_word = 8'hE0;
		16'h8479: out_word = 8'h04;
		16'h847A: out_word = 8'hE0;
		16'h847B: out_word = 8'h04;
		16'h847C: out_word = 8'hF3;
		16'h847D: out_word = 8'h04;
		16'h847E: out_word = 8'h01;
		16'h847F: out_word = 8'h05;
		16'h8480: out_word = 8'h12;
		16'h8481: out_word = 8'h05;
		16'h8482: out_word = 8'h23;
		16'h8483: out_word = 8'h05;
		16'h8484: out_word = 8'h31;
		16'h8485: out_word = 8'h05;
		16'h8486: out_word = 8'h42;
		16'h8487: out_word = 8'h05;
		16'h8488: out_word = 8'h4E;
		16'h8489: out_word = 8'h05;
		16'h848A: out_word = 8'h61;
		16'h848B: out_word = 8'h05;
		16'h848C: out_word = 8'h4D;
		16'h848D: out_word = 8'h45;
		16'h848E: out_word = 8'h52;
		16'h848F: out_word = 8'h47;
		16'h8490: out_word = 8'h45;
		16'h8491: out_word = 8'h20;
		16'h8492: out_word = 8'h65;
		16'h8493: out_word = 8'h72;
		16'h8494: out_word = 8'h72;
		16'h8495: out_word = 8'h6F;
		16'h8496: out_word = 8'hF2;
		16'h8497: out_word = 8'h57;
		16'h8498: out_word = 8'h72;
		16'h8499: out_word = 8'h6F;
		16'h849A: out_word = 8'h6E;
		16'h849B: out_word = 8'h67;
		16'h849C: out_word = 8'h20;
		16'h849D: out_word = 8'h66;
		16'h849E: out_word = 8'h69;
		16'h849F: out_word = 8'h6C;
		16'h84A0: out_word = 8'h65;
		16'h84A1: out_word = 8'h20;
		16'h84A2: out_word = 8'h74;
		16'h84A3: out_word = 8'h79;
		16'h84A4: out_word = 8'h70;
		16'h84A5: out_word = 8'hE5;
		16'h84A6: out_word = 8'h43;
		16'h84A7: out_word = 8'h4F;
		16'h84A8: out_word = 8'h44;
		16'h84A9: out_word = 8'h45;
		16'h84AA: out_word = 8'h20;
		16'h84AB: out_word = 8'h65;
		16'h84AC: out_word = 8'h72;
		16'h84AD: out_word = 8'h72;
		16'h84AE: out_word = 8'h6F;
		16'h84AF: out_word = 8'hF2;
		16'h84B0: out_word = 8'h54;
		16'h84B1: out_word = 8'h6F;
		16'h84B2: out_word = 8'h6F;
		16'h84B3: out_word = 8'h20;
		16'h84B4: out_word = 8'h6D;
		16'h84B5: out_word = 8'h61;
		16'h84B6: out_word = 8'h6E;
		16'h84B7: out_word = 8'h79;
		16'h84B8: out_word = 8'h20;
		16'h84B9: out_word = 8'h62;
		16'h84BA: out_word = 8'h72;
		16'h84BB: out_word = 8'h61;
		16'h84BC: out_word = 8'h63;
		16'h84BD: out_word = 8'h6B;
		16'h84BE: out_word = 8'h65;
		16'h84BF: out_word = 8'h74;
		16'h84C0: out_word = 8'hF3;
		16'h84C1: out_word = 8'h46;
		16'h84C2: out_word = 8'h69;
		16'h84C3: out_word = 8'h6C;
		16'h84C4: out_word = 8'h65;
		16'h84C5: out_word = 8'h20;
		16'h84C6: out_word = 8'h61;
		16'h84C7: out_word = 8'h6C;
		16'h84C8: out_word = 8'h72;
		16'h84C9: out_word = 8'h65;
		16'h84CA: out_word = 8'h61;
		16'h84CB: out_word = 8'h64;
		16'h84CC: out_word = 8'h79;
		16'h84CD: out_word = 8'h20;
		16'h84CE: out_word = 8'h65;
		16'h84CF: out_word = 8'h78;
		16'h84D0: out_word = 8'h69;
		16'h84D1: out_word = 8'h73;
		16'h84D2: out_word = 8'h74;
		16'h84D3: out_word = 8'hF3;
		16'h84D4: out_word = 8'h49;
		16'h84D5: out_word = 8'h6E;
		16'h84D6: out_word = 8'h76;
		16'h84D7: out_word = 8'h61;
		16'h84D8: out_word = 8'h6C;
		16'h84D9: out_word = 8'h69;
		16'h84DA: out_word = 8'h64;
		16'h84DB: out_word = 8'h20;
		16'h84DC: out_word = 8'h6E;
		16'h84DD: out_word = 8'h61;
		16'h84DE: out_word = 8'h6D;
		16'h84DF: out_word = 8'hE5;
		16'h84E0: out_word = 8'h46;
		16'h84E1: out_word = 8'h69;
		16'h84E2: out_word = 8'h6C;
		16'h84E3: out_word = 8'h65;
		16'h84E4: out_word = 8'h20;
		16'h84E5: out_word = 8'h64;
		16'h84E6: out_word = 8'h6F;
		16'h84E7: out_word = 8'h65;
		16'h84E8: out_word = 8'h73;
		16'h84E9: out_word = 8'h20;
		16'h84EA: out_word = 8'h6E;
		16'h84EB: out_word = 8'h6F;
		16'h84EC: out_word = 8'h74;
		16'h84ED: out_word = 8'h20;
		16'h84EE: out_word = 8'h65;
		16'h84EF: out_word = 8'h78;
		16'h84F0: out_word = 8'h69;
		16'h84F1: out_word = 8'h73;
		16'h84F2: out_word = 8'hF4;
		16'h84F3: out_word = 8'h49;
		16'h84F4: out_word = 8'h6E;
		16'h84F5: out_word = 8'h76;
		16'h84F6: out_word = 8'h61;
		16'h84F7: out_word = 8'h6C;
		16'h84F8: out_word = 8'h69;
		16'h84F9: out_word = 8'h64;
		16'h84FA: out_word = 8'h20;
		16'h84FB: out_word = 8'h64;
		16'h84FC: out_word = 8'h65;
		16'h84FD: out_word = 8'h76;
		16'h84FE: out_word = 8'h69;
		16'h84FF: out_word = 8'h63;
		16'h8500: out_word = 8'hE5;
		16'h8501: out_word = 8'h49;
		16'h8502: out_word = 8'h6E;
		16'h8503: out_word = 8'h76;
		16'h8504: out_word = 8'h61;
		16'h8505: out_word = 8'h6C;
		16'h8506: out_word = 8'h69;
		16'h8507: out_word = 8'h64;
		16'h8508: out_word = 8'h20;
		16'h8509: out_word = 8'h62;
		16'h850A: out_word = 8'h61;
		16'h850B: out_word = 8'h75;
		16'h850C: out_word = 8'h64;
		16'h850D: out_word = 8'h20;
		16'h850E: out_word = 8'h72;
		16'h850F: out_word = 8'h61;
		16'h8510: out_word = 8'h74;
		16'h8511: out_word = 8'hE5;
		16'h8512: out_word = 8'h49;
		16'h8513: out_word = 8'h6E;
		16'h8514: out_word = 8'h76;
		16'h8515: out_word = 8'h61;
		16'h8516: out_word = 8'h6C;
		16'h8517: out_word = 8'h69;
		16'h8518: out_word = 8'h64;
		16'h8519: out_word = 8'h20;
		16'h851A: out_word = 8'h6E;
		16'h851B: out_word = 8'h6F;
		16'h851C: out_word = 8'h74;
		16'h851D: out_word = 8'h65;
		16'h851E: out_word = 8'h20;
		16'h851F: out_word = 8'h6E;
		16'h8520: out_word = 8'h61;
		16'h8521: out_word = 8'h6D;
		16'h8522: out_word = 8'hE5;
		16'h8523: out_word = 8'h4E;
		16'h8524: out_word = 8'h75;
		16'h8525: out_word = 8'h6D;
		16'h8526: out_word = 8'h62;
		16'h8527: out_word = 8'h65;
		16'h8528: out_word = 8'h72;
		16'h8529: out_word = 8'h20;
		16'h852A: out_word = 8'h74;
		16'h852B: out_word = 8'h6F;
		16'h852C: out_word = 8'h6F;
		16'h852D: out_word = 8'h20;
		16'h852E: out_word = 8'h62;
		16'h852F: out_word = 8'h69;
		16'h8530: out_word = 8'hE7;
		16'h8531: out_word = 8'h4E;
		16'h8532: out_word = 8'h6F;
		16'h8533: out_word = 8'h74;
		16'h8534: out_word = 8'h65;
		16'h8535: out_word = 8'h20;
		16'h8536: out_word = 8'h6F;
		16'h8537: out_word = 8'h75;
		16'h8538: out_word = 8'h74;
		16'h8539: out_word = 8'h20;
		16'h853A: out_word = 8'h6F;
		16'h853B: out_word = 8'h66;
		16'h853C: out_word = 8'h20;
		16'h853D: out_word = 8'h72;
		16'h853E: out_word = 8'h61;
		16'h853F: out_word = 8'h6E;
		16'h8540: out_word = 8'h67;
		16'h8541: out_word = 8'hE5;
		16'h8542: out_word = 8'h4F;
		16'h8543: out_word = 8'h75;
		16'h8544: out_word = 8'h74;
		16'h8545: out_word = 8'h20;
		16'h8546: out_word = 8'h6F;
		16'h8547: out_word = 8'h66;
		16'h8548: out_word = 8'h20;
		16'h8549: out_word = 8'h72;
		16'h854A: out_word = 8'h61;
		16'h854B: out_word = 8'h6E;
		16'h854C: out_word = 8'h67;
		16'h854D: out_word = 8'hE5;
		16'h854E: out_word = 8'h54;
		16'h854F: out_word = 8'h6F;
		16'h8550: out_word = 8'h6F;
		16'h8551: out_word = 8'h20;
		16'h8552: out_word = 8'h6D;
		16'h8553: out_word = 8'h61;
		16'h8554: out_word = 8'h6E;
		16'h8555: out_word = 8'h79;
		16'h8556: out_word = 8'h20;
		16'h8557: out_word = 8'h74;
		16'h8558: out_word = 8'h69;
		16'h8559: out_word = 8'h65;
		16'h855A: out_word = 8'h64;
		16'h855B: out_word = 8'h20;
		16'h855C: out_word = 8'h6E;
		16'h855D: out_word = 8'h6F;
		16'h855E: out_word = 8'h74;
		16'h855F: out_word = 8'h65;
		16'h8560: out_word = 8'hF3;
		16'h8561: out_word = 8'h7F;
		16'h8562: out_word = 8'h20;
		16'h8563: out_word = 8'h31;
		16'h8564: out_word = 8'h39;
		16'h8565: out_word = 8'h38;
		16'h8566: out_word = 8'h36;
		16'h8567: out_word = 8'h20;
		16'h8568: out_word = 8'h53;
		16'h8569: out_word = 8'h69;
		16'h856A: out_word = 8'h6E;
		16'h856B: out_word = 8'h63;
		16'h856C: out_word = 8'h6C;
		16'h856D: out_word = 8'h61;
		16'h856E: out_word = 8'h69;
		16'h856F: out_word = 8'h72;
		16'h8570: out_word = 8'h20;
		16'h8571: out_word = 8'h52;
		16'h8572: out_word = 8'h65;
		16'h8573: out_word = 8'h73;
		16'h8574: out_word = 8'h65;
		16'h8575: out_word = 8'h61;
		16'h8576: out_word = 8'h72;
		16'h8577: out_word = 8'h63;
		16'h8578: out_word = 8'h68;
		16'h8579: out_word = 8'h20;
		16'h857A: out_word = 8'h4C;
		16'h857B: out_word = 8'h74;
		16'h857C: out_word = 8'hE4;
		16'h857D: out_word = 8'h1A;
		16'h857E: out_word = 8'hE6;
		16'h857F: out_word = 8'h7F;
		16'h8580: out_word = 8'hD5;
		16'h8581: out_word = 8'hD7;
		16'h8582: out_word = 8'hD1;
		16'h8583: out_word = 8'h1A;
		16'h8584: out_word = 8'h13;
		16'h8585: out_word = 8'h87;
		16'h8586: out_word = 8'h30;
		16'h8587: out_word = 8'hF5;
		16'h8588: out_word = 8'hC9;
		16'h8589: out_word = 8'hF4;
		16'h858A: out_word = 8'h09;
		16'h858B: out_word = 8'hA8;
		16'h858C: out_word = 8'h10;
		16'h858D: out_word = 8'h4B;
		16'h858E: out_word = 8'hF4;
		16'h858F: out_word = 8'h09;
		16'h8590: out_word = 8'hC4;
		16'h8591: out_word = 8'h15;
		16'h8592: out_word = 8'h53;
		16'h8593: out_word = 8'h81;
		16'h8594: out_word = 8'h0F;
		16'h8595: out_word = 8'hC4;
		16'h8596: out_word = 8'h15;
		16'h8597: out_word = 8'h52;
		16'h8598: out_word = 8'h34;
		16'h8599: out_word = 8'h5B;
		16'h859A: out_word = 8'h2F;
		16'h859B: out_word = 8'h5B;
		16'h859C: out_word = 8'h50;
		16'h859D: out_word = 8'h80;
		16'h859E: out_word = 8'h01;
		16'h859F: out_word = 8'h00;
		16'h85A0: out_word = 8'h06;
		16'h85A1: out_word = 8'h00;
		16'h85A2: out_word = 8'h0B;
		16'h85A3: out_word = 8'h00;
		16'h85A4: out_word = 8'h01;
		16'h85A5: out_word = 8'h00;
		16'h85A6: out_word = 8'h01;
		16'h85A7: out_word = 8'h00;
		16'h85A8: out_word = 8'h06;
		16'h85A9: out_word = 8'h00;
		16'h85AA: out_word = 8'h10;
		16'h85AB: out_word = 8'h00;
		16'h85AC: out_word = 8'hE1;
		16'h85AD: out_word = 8'h01;
		16'h85AE: out_word = 8'hFD;
		16'h85AF: out_word = 8'h7F;
		16'h85B0: out_word = 8'hAF;
		16'h85B1: out_word = 8'hF3;
		16'h85B2: out_word = 8'h32;
		16'h85B3: out_word = 8'h5C;
		16'h85B4: out_word = 8'h5B;
		16'h85B5: out_word = 8'hED;
		16'h85B6: out_word = 8'h79;
		16'h85B7: out_word = 8'hFB;
		16'h85B8: out_word = 8'hED;
		16'h85B9: out_word = 8'h7B;
		16'h85BA: out_word = 8'h3D;
		16'h85BB: out_word = 8'h5C;
		16'h85BC: out_word = 8'h7E;
		16'h85BD: out_word = 8'h32;
		16'h85BE: out_word = 8'h5E;
		16'h85BF: out_word = 8'h5B;
		16'h85C0: out_word = 8'h3C;
		16'h85C1: out_word = 8'hFE;
		16'h85C2: out_word = 8'h1E;
		16'h85C3: out_word = 8'h30;
		16'h85C4: out_word = 8'h03;
		16'h85C5: out_word = 8'hEF;
		16'h85C6: out_word = 8'h5D;
		16'h85C7: out_word = 8'h5B;
		16'h85C8: out_word = 8'h3D;
		16'h85C9: out_word = 8'hFD;
		16'h85CA: out_word = 8'h77;
		16'h85CB: out_word = 8'h00;
		16'h85CC: out_word = 8'h2A;
		16'h85CD: out_word = 8'h5D;
		16'h85CE: out_word = 8'h5C;
		16'h85CF: out_word = 8'h22;
		16'h85D0: out_word = 8'h5F;
		16'h85D1: out_word = 8'h5C;
		16'h85D2: out_word = 8'hEF;
		16'h85D3: out_word = 8'hC5;
		16'h85D4: out_word = 8'h16;
		16'h85D5: out_word = 8'hC9;
		16'h85D6: out_word = 8'h3E;
		16'h85D7: out_word = 8'h7F;
		16'h85D8: out_word = 8'hDB;
		16'h85D9: out_word = 8'hFE;
		16'h85DA: out_word = 8'h1F;
		16'h85DB: out_word = 8'hD8;
		16'h85DC: out_word = 8'h3E;
		16'h85DD: out_word = 8'hFE;
		16'h85DE: out_word = 8'hDB;
		16'h85DF: out_word = 8'hFE;
		16'h85E0: out_word = 8'h1F;
		16'h85E1: out_word = 8'hD8;
		16'h85E2: out_word = 8'hCD;
		16'h85E3: out_word = 8'hAC;
		16'h85E4: out_word = 8'h05;
		16'h85E5: out_word = 8'h14;
		16'h85E6: out_word = 8'hFB;
		16'h85E7: out_word = 8'h08;
		16'h85E8: out_word = 8'h11;
		16'h85E9: out_word = 8'h4A;
		16'h85EA: out_word = 8'h5B;
		16'h85EB: out_word = 8'hD5;
		16'h85EC: out_word = 8'hFD;
		16'h85ED: out_word = 8'hCB;
		16'h85EE: out_word = 8'h02;
		16'h85EF: out_word = 8'h9E;
		16'h85F0: out_word = 8'hE5;
		16'h85F1: out_word = 8'h2A;
		16'h85F2: out_word = 8'h3D;
		16'h85F3: out_word = 8'h5C;
		16'h85F4: out_word = 8'h5E;
		16'h85F5: out_word = 8'h23;
		16'h85F6: out_word = 8'h56;
		16'h85F7: out_word = 8'hA7;
		16'h85F8: out_word = 8'h21;
		16'h85F9: out_word = 8'h7F;
		16'h85FA: out_word = 8'h10;
		16'h85FB: out_word = 8'hED;
		16'h85FC: out_word = 8'h52;
		16'h85FD: out_word = 8'h20;
		16'h85FE: out_word = 8'h38;
		16'h85FF: out_word = 8'hE1;
		16'h8600: out_word = 8'hED;
		16'h8601: out_word = 8'h7B;
		16'h8602: out_word = 8'h3D;
		16'h8603: out_word = 8'h5C;
		16'h8604: out_word = 8'hD1;
		16'h8605: out_word = 8'hD1;
		16'h8606: out_word = 8'hED;
		16'h8607: out_word = 8'h53;
		16'h8608: out_word = 8'h3D;
		16'h8609: out_word = 8'h5C;
		16'h860A: out_word = 8'hE5;
		16'h860B: out_word = 8'h11;
		16'h860C: out_word = 8'h10;
		16'h860D: out_word = 8'h06;
		16'h860E: out_word = 8'hD5;
		16'h860F: out_word = 8'hE9;
		16'h8610: out_word = 8'h38;
		16'h8611: out_word = 8'h09;
		16'h8612: out_word = 8'h28;
		16'h8613: out_word = 8'h04;
		16'h8614: out_word = 8'hCD;
		16'h8615: out_word = 8'hAC;
		16'h8616: out_word = 8'h05;
		16'h8617: out_word = 8'h07;
		16'h8618: out_word = 8'hE1;
		16'h8619: out_word = 8'h18;
		16'h861A: out_word = 8'hEF;
		16'h861B: out_word = 8'hFE;
		16'h861C: out_word = 8'h0D;
		16'h861D: out_word = 8'h28;
		16'h861E: out_word = 8'h0E;
		16'h861F: out_word = 8'h2A;
		16'h8620: out_word = 8'h5A;
		16'h8621: out_word = 8'h5B;
		16'h8622: out_word = 8'hE5;
		16'h8623: out_word = 8'hEF;
		16'h8624: out_word = 8'h85;
		16'h8625: out_word = 8'h0F;
		16'h8626: out_word = 8'hE1;
		16'h8627: out_word = 8'h22;
		16'h8628: out_word = 8'h5A;
		16'h8629: out_word = 8'h5B;
		16'h862A: out_word = 8'hE1;
		16'h862B: out_word = 8'h18;
		16'h862C: out_word = 8'hDD;
		16'h862D: out_word = 8'hE1;
		16'h862E: out_word = 8'h3A;
		16'h862F: out_word = 8'h5C;
		16'h8630: out_word = 8'h5B;
		16'h8631: out_word = 8'hF6;
		16'h8632: out_word = 8'h10;
		16'h8633: out_word = 8'hF5;
		16'h8634: out_word = 8'hC3;
		16'h8635: out_word = 8'h4A;
		16'h8636: out_word = 8'h5B;
		16'h8637: out_word = 8'hE1;
		16'h8638: out_word = 8'h11;
		16'h8639: out_word = 8'h3D;
		16'h863A: out_word = 8'h06;
		16'h863B: out_word = 8'hD5;
		16'h863C: out_word = 8'hE9;
		16'h863D: out_word = 8'hD8;
		16'h863E: out_word = 8'hC8;
		16'h863F: out_word = 8'h18;
		16'h8640: out_word = 8'hD3;
		16'h8641: out_word = 8'hEF;
		16'h8642: out_word = 8'h18;
		16'h8643: out_word = 8'h00;
		16'h8644: out_word = 8'hEF;
		16'h8645: out_word = 8'h8C;
		16'h8646: out_word = 8'h1C;
		16'h8647: out_word = 8'hFD;
		16'h8648: out_word = 8'hCB;
		16'h8649: out_word = 8'h01;
		16'h864A: out_word = 8'h7E;
		16'h864B: out_word = 8'h28;
		16'h864C: out_word = 8'h14;
		16'h864D: out_word = 8'hEF;
		16'h864E: out_word = 8'hF1;
		16'h864F: out_word = 8'h2B;
		16'h8650: out_word = 8'h79;
		16'h8651: out_word = 8'h3D;
		16'h8652: out_word = 8'hB0;
		16'h8653: out_word = 8'h28;
		16'h8654: out_word = 8'h04;
		16'h8655: out_word = 8'hCD;
		16'h8656: out_word = 8'hAC;
		16'h8657: out_word = 8'h05;
		16'h8658: out_word = 8'h24;
		16'h8659: out_word = 8'h1A;
		16'h865A: out_word = 8'hE6;
		16'h865B: out_word = 8'hDF;
		16'h865C: out_word = 8'hFE;
		16'h865D: out_word = 8'h50;
		16'h865E: out_word = 8'hC2;
		16'h865F: out_word = 8'h12;
		16'h8660: out_word = 8'h19;
		16'h8661: out_word = 8'h2A;
		16'h8662: out_word = 8'h5D;
		16'h8663: out_word = 8'h5C;
		16'h8664: out_word = 8'h7E;
		16'h8665: out_word = 8'hFE;
		16'h8666: out_word = 8'h3B;
		16'h8667: out_word = 8'hC2;
		16'h8668: out_word = 8'h12;
		16'h8669: out_word = 8'h19;
		16'h866A: out_word = 8'hEF;
		16'h866B: out_word = 8'h20;
		16'h866C: out_word = 8'h00;
		16'h866D: out_word = 8'hEF;
		16'h866E: out_word = 8'h82;
		16'h866F: out_word = 8'h1C;
		16'h8670: out_word = 8'hFD;
		16'h8671: out_word = 8'hCB;
		16'h8672: out_word = 8'h01;
		16'h8673: out_word = 8'h7E;
		16'h8674: out_word = 8'h28;
		16'h8675: out_word = 8'h07;
		16'h8676: out_word = 8'hEF;
		16'h8677: out_word = 8'h99;
		16'h8678: out_word = 8'h1E;
		16'h8679: out_word = 8'hED;
		16'h867A: out_word = 8'h43;
		16'h867B: out_word = 8'h71;
		16'h867C: out_word = 8'h5B;
		16'h867D: out_word = 8'hEF;
		16'h867E: out_word = 8'h18;
		16'h867F: out_word = 8'h00;
		16'h8680: out_word = 8'hFE;
		16'h8681: out_word = 8'h0D;
		16'h8682: out_word = 8'h28;
		16'h8683: out_word = 8'h05;
		16'h8684: out_word = 8'hFE;
		16'h8685: out_word = 8'h3A;
		16'h8686: out_word = 8'hC2;
		16'h8687: out_word = 8'h12;
		16'h8688: out_word = 8'h19;
		16'h8689: out_word = 8'hCD;
		16'h868A: out_word = 8'hA1;
		16'h868B: out_word = 8'h18;
		16'h868C: out_word = 8'hED;
		16'h868D: out_word = 8'h4B;
		16'h868E: out_word = 8'h71;
		16'h868F: out_word = 8'h5B;
		16'h8690: out_word = 8'h78;
		16'h8691: out_word = 8'hB1;
		16'h8692: out_word = 8'h20;
		16'h8693: out_word = 8'h04;
		16'h8694: out_word = 8'hCD;
		16'h8695: out_word = 8'hAC;
		16'h8696: out_word = 8'h05;
		16'h8697: out_word = 8'h25;
		16'h8698: out_word = 8'h21;
		16'h8699: out_word = 8'hB8;
		16'h869A: out_word = 8'h06;
		16'h869B: out_word = 8'h5E;
		16'h869C: out_word = 8'h23;
		16'h869D: out_word = 8'h56;
		16'h869E: out_word = 8'h23;
		16'h869F: out_word = 8'hEB;
		16'h86A0: out_word = 8'h7C;
		16'h86A1: out_word = 8'hFE;
		16'h86A2: out_word = 8'h25;
		16'h86A3: out_word = 8'h30;
		16'h86A4: out_word = 8'h0A;
		16'h86A5: out_word = 8'hA7;
		16'h86A6: out_word = 8'hED;
		16'h86A7: out_word = 8'h42;
		16'h86A8: out_word = 8'h30;
		16'h86A9: out_word = 8'h05;
		16'h86AA: out_word = 8'hEB;
		16'h86AB: out_word = 8'h23;
		16'h86AC: out_word = 8'h23;
		16'h86AD: out_word = 8'h18;
		16'h86AE: out_word = 8'hEC;
		16'h86AF: out_word = 8'hEB;
		16'h86B0: out_word = 8'h5E;
		16'h86B1: out_word = 8'h23;
		16'h86B2: out_word = 8'h56;
		16'h86B3: out_word = 8'hED;
		16'h86B4: out_word = 8'h53;
		16'h86B5: out_word = 8'h5F;
		16'h86B6: out_word = 8'h5B;
		16'h86B7: out_word = 8'hC9;
		16'h86B8: out_word = 8'h32;
		16'h86B9: out_word = 8'h00;
		16'h86BA: out_word = 8'hA5;
		16'h86BB: out_word = 8'h0A;
		16'h86BC: out_word = 8'h6E;
		16'h86BD: out_word = 8'h00;
		16'h86BE: out_word = 8'hD4;
		16'h86BF: out_word = 8'h04;
		16'h86C0: out_word = 8'h2C;
		16'h86C1: out_word = 8'h01;
		16'h86C2: out_word = 8'hC3;
		16'h86C3: out_word = 8'h01;
		16'h86C4: out_word = 8'h58;
		16'h86C5: out_word = 8'h02;
		16'h86C6: out_word = 8'hE0;
		16'h86C7: out_word = 8'h00;
		16'h86C8: out_word = 8'hB0;
		16'h86C9: out_word = 8'h04;
		16'h86CA: out_word = 8'h6E;
		16'h86CB: out_word = 8'h00;
		16'h86CC: out_word = 8'h60;
		16'h86CD: out_word = 8'h09;
		16'h86CE: out_word = 8'h36;
		16'h86CF: out_word = 8'h00;
		16'h86D0: out_word = 8'hC0;
		16'h86D1: out_word = 8'h12;
		16'h86D2: out_word = 8'h19;
		16'h86D3: out_word = 8'h00;
		16'h86D4: out_word = 8'h80;
		16'h86D5: out_word = 8'h25;
		16'h86D6: out_word = 8'h0B;
		16'h86D7: out_word = 8'h00;
		16'h86D8: out_word = 8'h21;
		16'h86D9: out_word = 8'h61;
		16'h86DA: out_word = 8'h5B;
		16'h86DB: out_word = 8'h7E;
		16'h86DC: out_word = 8'hA7;
		16'h86DD: out_word = 8'h28;
		16'h86DE: out_word = 8'h06;
		16'h86DF: out_word = 8'h36;
		16'h86E0: out_word = 8'h00;
		16'h86E1: out_word = 8'h23;
		16'h86E2: out_word = 8'h7E;
		16'h86E3: out_word = 8'h37;
		16'h86E4: out_word = 8'hC9;
		16'h86E5: out_word = 8'hCD;
		16'h86E6: out_word = 8'hD6;
		16'h86E7: out_word = 8'h05;
		16'h86E8: out_word = 8'hF3;
		16'h86E9: out_word = 8'hD9;
		16'h86EA: out_word = 8'hED;
		16'h86EB: out_word = 8'h5B;
		16'h86EC: out_word = 8'h5F;
		16'h86ED: out_word = 8'h5B;
		16'h86EE: out_word = 8'h2A;
		16'h86EF: out_word = 8'h5F;
		16'h86F0: out_word = 8'h5B;
		16'h86F1: out_word = 8'hCB;
		16'h86F2: out_word = 8'h3C;
		16'h86F3: out_word = 8'hCB;
		16'h86F4: out_word = 8'h1D;
		16'h86F5: out_word = 8'hB7;
		16'h86F6: out_word = 8'h06;
		16'h86F7: out_word = 8'hFA;
		16'h86F8: out_word = 8'hD9;
		16'h86F9: out_word = 8'h0E;
		16'h86FA: out_word = 8'hFD;
		16'h86FB: out_word = 8'h16;
		16'h86FC: out_word = 8'hFF;
		16'h86FD: out_word = 8'h1E;
		16'h86FE: out_word = 8'hBF;
		16'h86FF: out_word = 8'h42;
		16'h8700: out_word = 8'h3E;
		16'h8701: out_word = 8'h0E;
		16'h8702: out_word = 8'hED;
		16'h8703: out_word = 8'h79;
		16'h8704: out_word = 8'hED;
		16'h8705: out_word = 8'h78;
		16'h8706: out_word = 8'hF6;
		16'h8707: out_word = 8'hF0;
		16'h8708: out_word = 8'hE6;
		16'h8709: out_word = 8'hFB;
		16'h870A: out_word = 8'h43;
		16'h870B: out_word = 8'hED;
		16'h870C: out_word = 8'h79;
		16'h870D: out_word = 8'h67;
		16'h870E: out_word = 8'h42;
		16'h870F: out_word = 8'hED;
		16'h8710: out_word = 8'h78;
		16'h8711: out_word = 8'hE6;
		16'h8712: out_word = 8'h80;
		16'h8713: out_word = 8'h28;
		16'h8714: out_word = 8'h09;
		16'h8715: out_word = 8'hD9;
		16'h8716: out_word = 8'h05;
		16'h8717: out_word = 8'hD9;
		16'h8718: out_word = 8'h20;
		16'h8719: out_word = 8'hF4;
		16'h871A: out_word = 8'hAF;
		16'h871B: out_word = 8'hF5;
		16'h871C: out_word = 8'h18;
		16'h871D: out_word = 8'h39;
		16'h871E: out_word = 8'hED;
		16'h871F: out_word = 8'h78;
		16'h8720: out_word = 8'hE6;
		16'h8721: out_word = 8'h80;
		16'h8722: out_word = 8'h20;
		16'h8723: out_word = 8'hF1;
		16'h8724: out_word = 8'hED;
		16'h8725: out_word = 8'h78;
		16'h8726: out_word = 8'hE6;
		16'h8727: out_word = 8'h80;
		16'h8728: out_word = 8'h20;
		16'h8729: out_word = 8'hEB;
		16'h872A: out_word = 8'hD9;
		16'h872B: out_word = 8'h01;
		16'h872C: out_word = 8'hFD;
		16'h872D: out_word = 8'hFF;
		16'h872E: out_word = 8'h3E;
		16'h872F: out_word = 8'h80;
		16'h8730: out_word = 8'h08;
		16'h8731: out_word = 8'h19;
		16'h8732: out_word = 8'h00;
		16'h8733: out_word = 8'h00;
		16'h8734: out_word = 8'h00;
		16'h8735: out_word = 8'h00;
		16'h8736: out_word = 8'h2B;
		16'h8737: out_word = 8'h7C;
		16'h8738: out_word = 8'hB5;
		16'h8739: out_word = 8'h20;
		16'h873A: out_word = 8'hFB;
		16'h873B: out_word = 8'hED;
		16'h873C: out_word = 8'h78;
		16'h873D: out_word = 8'hE6;
		16'h873E: out_word = 8'h80;
		16'h873F: out_word = 8'hCA;
		16'h8740: out_word = 8'h4B;
		16'h8741: out_word = 8'h07;
		16'h8742: out_word = 8'h08;
		16'h8743: out_word = 8'h37;
		16'h8744: out_word = 8'h1F;
		16'h8745: out_word = 8'h38;
		16'h8746: out_word = 8'h0D;
		16'h8747: out_word = 8'h08;
		16'h8748: out_word = 8'hC3;
		16'h8749: out_word = 8'h31;
		16'h874A: out_word = 8'h07;
		16'h874B: out_word = 8'h08;
		16'h874C: out_word = 8'hB7;
		16'h874D: out_word = 8'h1F;
		16'h874E: out_word = 8'h38;
		16'h874F: out_word = 8'h04;
		16'h8750: out_word = 8'h08;
		16'h8751: out_word = 8'hC3;
		16'h8752: out_word = 8'h31;
		16'h8753: out_word = 8'h07;
		16'h8754: out_word = 8'h37;
		16'h8755: out_word = 8'hF5;
		16'h8756: out_word = 8'hD9;
		16'h8757: out_word = 8'h7C;
		16'h8758: out_word = 8'hF6;
		16'h8759: out_word = 8'h04;
		16'h875A: out_word = 8'h43;
		16'h875B: out_word = 8'hED;
		16'h875C: out_word = 8'h79;
		16'h875D: out_word = 8'hD9;
		16'h875E: out_word = 8'h62;
		16'h875F: out_word = 8'h6B;
		16'h8760: out_word = 8'h01;
		16'h8761: out_word = 8'h07;
		16'h8762: out_word = 8'h00;
		16'h8763: out_word = 8'hB7;
		16'h8764: out_word = 8'hED;
		16'h8765: out_word = 8'h42;
		16'h8766: out_word = 8'h2B;
		16'h8767: out_word = 8'h7C;
		16'h8768: out_word = 8'hB5;
		16'h8769: out_word = 8'h20;
		16'h876A: out_word = 8'hFB;
		16'h876B: out_word = 8'h01;
		16'h876C: out_word = 8'hFD;
		16'h876D: out_word = 8'hFF;
		16'h876E: out_word = 8'h19;
		16'h876F: out_word = 8'h19;
		16'h8770: out_word = 8'h19;
		16'h8771: out_word = 8'hED;
		16'h8772: out_word = 8'h78;
		16'h8773: out_word = 8'hE6;
		16'h8774: out_word = 8'h80;
		16'h8775: out_word = 8'h28;
		16'h8776: out_word = 8'h08;
		16'h8777: out_word = 8'h2B;
		16'h8778: out_word = 8'h7C;
		16'h8779: out_word = 8'hB5;
		16'h877A: out_word = 8'h20;
		16'h877B: out_word = 8'hF5;
		16'h877C: out_word = 8'hF1;
		16'h877D: out_word = 8'hFB;
		16'h877E: out_word = 8'hC9;
		16'h877F: out_word = 8'hED;
		16'h8780: out_word = 8'h78;
		16'h8781: out_word = 8'hE6;
		16'h8782: out_word = 8'h80;
		16'h8783: out_word = 8'h20;
		16'h8784: out_word = 8'hEC;
		16'h8785: out_word = 8'hED;
		16'h8786: out_word = 8'h78;
		16'h8787: out_word = 8'hE6;
		16'h8788: out_word = 8'h80;
		16'h8789: out_word = 8'h20;
		16'h878A: out_word = 8'hE6;
		16'h878B: out_word = 8'h62;
		16'h878C: out_word = 8'h6B;
		16'h878D: out_word = 8'h01;
		16'h878E: out_word = 8'h02;
		16'h878F: out_word = 8'h00;
		16'h8790: out_word = 8'hCB;
		16'h8791: out_word = 8'h3C;
		16'h8792: out_word = 8'hCB;
		16'h8793: out_word = 8'h1D;
		16'h8794: out_word = 8'hB7;
		16'h8795: out_word = 8'hED;
		16'h8796: out_word = 8'h42;
		16'h8797: out_word = 8'h01;
		16'h8798: out_word = 8'hFD;
		16'h8799: out_word = 8'hFF;
		16'h879A: out_word = 8'h3E;
		16'h879B: out_word = 8'h80;
		16'h879C: out_word = 8'h08;
		16'h879D: out_word = 8'h00;
		16'h879E: out_word = 8'h00;
		16'h879F: out_word = 8'h00;
		16'h87A0: out_word = 8'h00;
		16'h87A1: out_word = 8'h19;
		16'h87A2: out_word = 8'h2B;
		16'h87A3: out_word = 8'h7C;
		16'h87A4: out_word = 8'hB5;
		16'h87A5: out_word = 8'h20;
		16'h87A6: out_word = 8'hFB;
		16'h87A7: out_word = 8'hED;
		16'h87A8: out_word = 8'h78;
		16'h87A9: out_word = 8'hE6;
		16'h87AA: out_word = 8'h80;
		16'h87AB: out_word = 8'hCA;
		16'h87AC: out_word = 8'hB7;
		16'h87AD: out_word = 8'h07;
		16'h87AE: out_word = 8'h08;
		16'h87AF: out_word = 8'h37;
		16'h87B0: out_word = 8'h1F;
		16'h87B1: out_word = 8'h38;
		16'h87B2: out_word = 8'h0D;
		16'h87B3: out_word = 8'h08;
		16'h87B4: out_word = 8'hC3;
		16'h87B5: out_word = 8'h9D;
		16'h87B6: out_word = 8'h07;
		16'h87B7: out_word = 8'h08;
		16'h87B8: out_word = 8'hB7;
		16'h87B9: out_word = 8'h1F;
		16'h87BA: out_word = 8'h38;
		16'h87BB: out_word = 8'h04;
		16'h87BC: out_word = 8'h08;
		16'h87BD: out_word = 8'hC3;
		16'h87BE: out_word = 8'h9D;
		16'h87BF: out_word = 8'h07;
		16'h87C0: out_word = 8'h21;
		16'h87C1: out_word = 8'h61;
		16'h87C2: out_word = 8'h5B;
		16'h87C3: out_word = 8'h36;
		16'h87C4: out_word = 8'h01;
		16'h87C5: out_word = 8'h23;
		16'h87C6: out_word = 8'h77;
		16'h87C7: out_word = 8'hF1;
		16'h87C8: out_word = 8'hFB;
		16'h87C9: out_word = 8'hC9;
		16'h87CA: out_word = 8'hF5;
		16'h87CB: out_word = 8'h3A;
		16'h87CC: out_word = 8'h65;
		16'h87CD: out_word = 8'h5B;
		16'h87CE: out_word = 8'hB7;
		16'h87CF: out_word = 8'h28;
		16'h87D0: out_word = 8'h0F;
		16'h87D1: out_word = 8'h3D;
		16'h87D2: out_word = 8'h32;
		16'h87D3: out_word = 8'h65;
		16'h87D4: out_word = 8'h5B;
		16'h87D5: out_word = 8'h20;
		16'h87D6: out_word = 8'h04;
		16'h87D7: out_word = 8'hF1;
		16'h87D8: out_word = 8'hC3;
		16'h87D9: out_word = 8'h72;
		16'h87DA: out_word = 8'h08;
		16'h87DB: out_word = 8'hF1;
		16'h87DC: out_word = 8'h32;
		16'h87DD: out_word = 8'h0F;
		16'h87DE: out_word = 8'h5C;
		16'h87DF: out_word = 8'hC9;
		16'h87E0: out_word = 8'hF1;
		16'h87E1: out_word = 8'hFE;
		16'h87E2: out_word = 8'hA3;
		16'h87E3: out_word = 8'h38;
		16'h87E4: out_word = 8'h0D;
		16'h87E5: out_word = 8'h2A;
		16'h87E6: out_word = 8'h5A;
		16'h87E7: out_word = 8'h5B;
		16'h87E8: out_word = 8'hE5;
		16'h87E9: out_word = 8'hEF;
		16'h87EA: out_word = 8'h52;
		16'h87EB: out_word = 8'h0B;
		16'h87EC: out_word = 8'hE1;
		16'h87ED: out_word = 8'h22;
		16'h87EE: out_word = 8'h5A;
		16'h87EF: out_word = 8'h5B;
		16'h87F0: out_word = 8'h37;
		16'h87F1: out_word = 8'hC9;
		16'h87F2: out_word = 8'h21;
		16'h87F3: out_word = 8'h3B;
		16'h87F4: out_word = 8'h5C;
		16'h87F5: out_word = 8'hCB;
		16'h87F6: out_word = 8'h86;
		16'h87F7: out_word = 8'hFE;
		16'h87F8: out_word = 8'h20;
		16'h87F9: out_word = 8'h20;
		16'h87FA: out_word = 8'h02;
		16'h87FB: out_word = 8'hCB;
		16'h87FC: out_word = 8'hC6;
		16'h87FD: out_word = 8'hFE;
		16'h87FE: out_word = 8'h7F;
		16'h87FF: out_word = 8'h38;
		16'h8800: out_word = 8'h02;
		16'h8801: out_word = 8'h3E;
		16'h8802: out_word = 8'h3F;
		16'h8803: out_word = 8'hFE;
		16'h8804: out_word = 8'h20;
		16'h8805: out_word = 8'h38;
		16'h8806: out_word = 8'h17;
		16'h8807: out_word = 8'hF5;
		16'h8808: out_word = 8'h21;
		16'h8809: out_word = 8'h63;
		16'h880A: out_word = 8'h5B;
		16'h880B: out_word = 8'h34;
		16'h880C: out_word = 8'h3A;
		16'h880D: out_word = 8'h64;
		16'h880E: out_word = 8'h5B;
		16'h880F: out_word = 8'hBE;
		16'h8810: out_word = 8'h30;
		16'h8811: out_word = 8'h08;
		16'h8812: out_word = 8'hCD;
		16'h8813: out_word = 8'h22;
		16'h8814: out_word = 8'h08;
		16'h8815: out_word = 8'h3E;
		16'h8816: out_word = 8'h01;
		16'h8817: out_word = 8'h32;
		16'h8818: out_word = 8'h63;
		16'h8819: out_word = 8'h5B;
		16'h881A: out_word = 8'hF1;
		16'h881B: out_word = 8'hC3;
		16'h881C: out_word = 8'hA3;
		16'h881D: out_word = 8'h08;
		16'h881E: out_word = 8'hFE;
		16'h881F: out_word = 8'h0D;
		16'h8820: out_word = 8'h20;
		16'h8821: out_word = 8'h0E;
		16'h8822: out_word = 8'hAF;
		16'h8823: out_word = 8'h32;
		16'h8824: out_word = 8'h63;
		16'h8825: out_word = 8'h5B;
		16'h8826: out_word = 8'h3E;
		16'h8827: out_word = 8'h0D;
		16'h8828: out_word = 8'hCD;
		16'h8829: out_word = 8'hA3;
		16'h882A: out_word = 8'h08;
		16'h882B: out_word = 8'h3E;
		16'h882C: out_word = 8'h0A;
		16'h882D: out_word = 8'hC3;
		16'h882E: out_word = 8'hA3;
		16'h882F: out_word = 8'h08;
		16'h8830: out_word = 8'hFE;
		16'h8831: out_word = 8'h06;
		16'h8832: out_word = 8'h20;
		16'h8833: out_word = 8'h1F;
		16'h8834: out_word = 8'hED;
		16'h8835: out_word = 8'h4B;
		16'h8836: out_word = 8'h63;
		16'h8837: out_word = 8'h5B;
		16'h8838: out_word = 8'h1E;
		16'h8839: out_word = 8'h00;
		16'h883A: out_word = 8'h1C;
		16'h883B: out_word = 8'h0C;
		16'h883C: out_word = 8'h79;
		16'h883D: out_word = 8'hB8;
		16'h883E: out_word = 8'h28;
		16'h883F: out_word = 8'h08;
		16'h8840: out_word = 8'hD6;
		16'h8841: out_word = 8'h08;
		16'h8842: out_word = 8'h28;
		16'h8843: out_word = 8'h04;
		16'h8844: out_word = 8'h30;
		16'h8845: out_word = 8'hFA;
		16'h8846: out_word = 8'h18;
		16'h8847: out_word = 8'hF2;
		16'h8848: out_word = 8'hD5;
		16'h8849: out_word = 8'h3E;
		16'h884A: out_word = 8'h20;
		16'h884B: out_word = 8'hCD;
		16'h884C: out_word = 8'hCA;
		16'h884D: out_word = 8'h07;
		16'h884E: out_word = 8'hD1;
		16'h884F: out_word = 8'h1D;
		16'h8850: out_word = 8'hC8;
		16'h8851: out_word = 8'h18;
		16'h8852: out_word = 8'hF5;
		16'h8853: out_word = 8'hFE;
		16'h8854: out_word = 8'h16;
		16'h8855: out_word = 8'h28;
		16'h8856: out_word = 8'h09;
		16'h8857: out_word = 8'hFE;
		16'h8858: out_word = 8'h17;
		16'h8859: out_word = 8'h28;
		16'h885A: out_word = 8'h05;
		16'h885B: out_word = 8'hFE;
		16'h885C: out_word = 8'h10;
		16'h885D: out_word = 8'hD8;
		16'h885E: out_word = 8'h18;
		16'h885F: out_word = 8'h09;
		16'h8860: out_word = 8'h32;
		16'h8861: out_word = 8'h0E;
		16'h8862: out_word = 8'h5C;
		16'h8863: out_word = 8'h3E;
		16'h8864: out_word = 8'h02;
		16'h8865: out_word = 8'h32;
		16'h8866: out_word = 8'h65;
		16'h8867: out_word = 8'h5B;
		16'h8868: out_word = 8'hC9;
		16'h8869: out_word = 8'h32;
		16'h886A: out_word = 8'h0E;
		16'h886B: out_word = 8'h5C;
		16'h886C: out_word = 8'h3E;
		16'h886D: out_word = 8'h02;
		16'h886E: out_word = 8'h32;
		16'h886F: out_word = 8'h65;
		16'h8870: out_word = 8'h5B;
		16'h8871: out_word = 8'hC9;
		16'h8872: out_word = 8'h57;
		16'h8873: out_word = 8'h3A;
		16'h8874: out_word = 8'h0E;
		16'h8875: out_word = 8'h5C;
		16'h8876: out_word = 8'hFE;
		16'h8877: out_word = 8'h16;
		16'h8878: out_word = 8'h28;
		16'h8879: out_word = 8'h08;
		16'h887A: out_word = 8'hFE;
		16'h887B: out_word = 8'h17;
		16'h887C: out_word = 8'h3F;
		16'h887D: out_word = 8'hC0;
		16'h887E: out_word = 8'h3A;
		16'h887F: out_word = 8'h0F;
		16'h8880: out_word = 8'h5C;
		16'h8881: out_word = 8'h57;
		16'h8882: out_word = 8'h3A;
		16'h8883: out_word = 8'h64;
		16'h8884: out_word = 8'h5B;
		16'h8885: out_word = 8'hBA;
		16'h8886: out_word = 8'h28;
		16'h8887: out_word = 8'h02;
		16'h8888: out_word = 8'h30;
		16'h8889: out_word = 8'h06;
		16'h888A: out_word = 8'h47;
		16'h888B: out_word = 8'h7A;
		16'h888C: out_word = 8'h90;
		16'h888D: out_word = 8'h57;
		16'h888E: out_word = 8'h18;
		16'h888F: out_word = 8'hF2;
		16'h8890: out_word = 8'h7A;
		16'h8891: out_word = 8'hB7;
		16'h8892: out_word = 8'hCA;
		16'h8893: out_word = 8'h22;
		16'h8894: out_word = 8'h08;
		16'h8895: out_word = 8'h3A;
		16'h8896: out_word = 8'h63;
		16'h8897: out_word = 8'h5B;
		16'h8898: out_word = 8'hBA;
		16'h8899: out_word = 8'hC8;
		16'h889A: out_word = 8'hD5;
		16'h889B: out_word = 8'h3E;
		16'h889C: out_word = 8'h20;
		16'h889D: out_word = 8'hCD;
		16'h889E: out_word = 8'hCA;
		16'h889F: out_word = 8'h07;
		16'h88A0: out_word = 8'hD1;
		16'h88A1: out_word = 8'h18;
		16'h88A2: out_word = 8'hF2;
		16'h88A3: out_word = 8'hF5;
		16'h88A4: out_word = 8'h0E;
		16'h88A5: out_word = 8'hFD;
		16'h88A6: out_word = 8'h16;
		16'h88A7: out_word = 8'hFF;
		16'h88A8: out_word = 8'h1E;
		16'h88A9: out_word = 8'hBF;
		16'h88AA: out_word = 8'h42;
		16'h88AB: out_word = 8'h3E;
		16'h88AC: out_word = 8'h0E;
		16'h88AD: out_word = 8'hED;
		16'h88AE: out_word = 8'h79;
		16'h88AF: out_word = 8'hCD;
		16'h88B0: out_word = 8'hD6;
		16'h88B1: out_word = 8'h05;
		16'h88B2: out_word = 8'hED;
		16'h88B3: out_word = 8'h78;
		16'h88B4: out_word = 8'hE6;
		16'h88B5: out_word = 8'h40;
		16'h88B6: out_word = 8'h20;
		16'h88B7: out_word = 8'hF7;
		16'h88B8: out_word = 8'h2A;
		16'h88B9: out_word = 8'h5F;
		16'h88BA: out_word = 8'h5B;
		16'h88BB: out_word = 8'h11;
		16'h88BC: out_word = 8'h02;
		16'h88BD: out_word = 8'h00;
		16'h88BE: out_word = 8'hB7;
		16'h88BF: out_word = 8'hED;
		16'h88C0: out_word = 8'h52;
		16'h88C1: out_word = 8'hEB;
		16'h88C2: out_word = 8'hF1;
		16'h88C3: out_word = 8'h2F;
		16'h88C4: out_word = 8'h37;
		16'h88C5: out_word = 8'h06;
		16'h88C6: out_word = 8'h0B;
		16'h88C7: out_word = 8'hF3;
		16'h88C8: out_word = 8'hC5;
		16'h88C9: out_word = 8'hF5;
		16'h88CA: out_word = 8'h3E;
		16'h88CB: out_word = 8'hFE;
		16'h88CC: out_word = 8'h62;
		16'h88CD: out_word = 8'h6B;
		16'h88CE: out_word = 8'h01;
		16'h88CF: out_word = 8'hFD;
		16'h88D0: out_word = 8'hBF;
		16'h88D1: out_word = 8'hD2;
		16'h88D2: out_word = 8'hDA;
		16'h88D3: out_word = 8'h08;
		16'h88D4: out_word = 8'hE6;
		16'h88D5: out_word = 8'hF7;
		16'h88D6: out_word = 8'hED;
		16'h88D7: out_word = 8'h79;
		16'h88D8: out_word = 8'h18;
		16'h88D9: out_word = 8'h06;
		16'h88DA: out_word = 8'hF6;
		16'h88DB: out_word = 8'h08;
		16'h88DC: out_word = 8'hED;
		16'h88DD: out_word = 8'h79;
		16'h88DE: out_word = 8'h18;
		16'h88DF: out_word = 8'h00;
		16'h88E0: out_word = 8'h2B;
		16'h88E1: out_word = 8'h7C;
		16'h88E2: out_word = 8'hB5;
		16'h88E3: out_word = 8'h20;
		16'h88E4: out_word = 8'hFB;
		16'h88E5: out_word = 8'h00;
		16'h88E6: out_word = 8'h00;
		16'h88E7: out_word = 8'h00;
		16'h88E8: out_word = 8'hF1;
		16'h88E9: out_word = 8'hC1;
		16'h88EA: out_word = 8'hB7;
		16'h88EB: out_word = 8'h1F;
		16'h88EC: out_word = 8'h10;
		16'h88ED: out_word = 8'hDA;
		16'h88EE: out_word = 8'hFB;
		16'h88EF: out_word = 8'hC9;
		16'h88F0: out_word = 8'h21;
		16'h88F1: out_word = 8'h72;
		16'h88F2: out_word = 8'h5B;
		16'h88F3: out_word = 8'h36;
		16'h88F4: out_word = 8'h2B;
		16'h88F5: out_word = 8'h21;
		16'h88F6: out_word = 8'h79;
		16'h88F7: out_word = 8'h09;
		16'h88F8: out_word = 8'hCD;
		16'h88F9: out_word = 8'h5F;
		16'h88FA: out_word = 8'h09;
		16'h88FB: out_word = 8'hCD;
		16'h88FC: out_word = 8'h15;
		16'h88FD: out_word = 8'h09;
		16'h88FE: out_word = 8'h21;
		16'h88FF: out_word = 8'h80;
		16'h8900: out_word = 8'h09;
		16'h8901: out_word = 8'hCD;
		16'h8902: out_word = 8'h5F;
		16'h8903: out_word = 8'h09;
		16'h8904: out_word = 8'h21;
		16'h8905: out_word = 8'h72;
		16'h8906: out_word = 8'h5B;
		16'h8907: out_word = 8'hAF;
		16'h8908: out_word = 8'hBE;
		16'h8909: out_word = 8'h28;
		16'h890A: out_word = 8'h03;
		16'h890B: out_word = 8'h35;
		16'h890C: out_word = 8'h18;
		16'h890D: out_word = 8'hE7;
		16'h890E: out_word = 8'h21;
		16'h890F: out_word = 8'h82;
		16'h8910: out_word = 8'h09;
		16'h8911: out_word = 8'hCD;
		16'h8912: out_word = 8'h5F;
		16'h8913: out_word = 8'h09;
		16'h8914: out_word = 8'hC9;
		16'h8915: out_word = 8'h21;
		16'h8916: out_word = 8'h71;
		16'h8917: out_word = 8'h5B;
		16'h8918: out_word = 8'h36;
		16'h8919: out_word = 8'hFF;
		16'h891A: out_word = 8'hCD;
		16'h891B: out_word = 8'h26;
		16'h891C: out_word = 8'h09;
		16'h891D: out_word = 8'h21;
		16'h891E: out_word = 8'h71;
		16'h891F: out_word = 8'h5B;
		16'h8920: out_word = 8'hAF;
		16'h8921: out_word = 8'hBE;
		16'h8922: out_word = 8'hC8;
		16'h8923: out_word = 8'h35;
		16'h8924: out_word = 8'h18;
		16'h8925: out_word = 8'hF4;
		16'h8926: out_word = 8'h11;
		16'h8927: out_word = 8'h00;
		16'h8928: out_word = 8'hC0;
		16'h8929: out_word = 8'hED;
		16'h892A: out_word = 8'h4B;
		16'h892B: out_word = 8'h71;
		16'h892C: out_word = 8'h5B;
		16'h892D: out_word = 8'h37;
		16'h892E: out_word = 8'hCB;
		16'h892F: out_word = 8'h10;
		16'h8930: out_word = 8'h37;
		16'h8931: out_word = 8'hCB;
		16'h8932: out_word = 8'h10;
		16'h8933: out_word = 8'h79;
		16'h8934: out_word = 8'h2F;
		16'h8935: out_word = 8'h4F;
		16'h8936: out_word = 8'hAF;
		16'h8937: out_word = 8'hF5;
		16'h8938: out_word = 8'hD5;
		16'h8939: out_word = 8'hC5;
		16'h893A: out_word = 8'hCD;
		16'h893B: out_word = 8'h6D;
		16'h893C: out_word = 8'h09;
		16'h893D: out_word = 8'hC1;
		16'h893E: out_word = 8'hD1;
		16'h893F: out_word = 8'h1E;
		16'h8940: out_word = 8'h00;
		16'h8941: out_word = 8'h28;
		16'h8942: out_word = 8'h01;
		16'h8943: out_word = 8'h5A;
		16'h8944: out_word = 8'hF1;
		16'h8945: out_word = 8'hB3;
		16'h8946: out_word = 8'hF5;
		16'h8947: out_word = 8'h05;
		16'h8948: out_word = 8'hCB;
		16'h8949: out_word = 8'h3A;
		16'h894A: out_word = 8'hCB;
		16'h894B: out_word = 8'h3A;
		16'h894C: out_word = 8'hD5;
		16'h894D: out_word = 8'hC5;
		16'h894E: out_word = 8'h30;
		16'h894F: out_word = 8'hEA;
		16'h8950: out_word = 8'hC1;
		16'h8951: out_word = 8'hD1;
		16'h8952: out_word = 8'hF1;
		16'h8953: out_word = 8'h06;
		16'h8954: out_word = 8'h03;
		16'h8955: out_word = 8'hC5;
		16'h8956: out_word = 8'hF5;
		16'h8957: out_word = 8'hCD;
		16'h8958: out_word = 8'hA3;
		16'h8959: out_word = 8'h08;
		16'h895A: out_word = 8'hF1;
		16'h895B: out_word = 8'hC1;
		16'h895C: out_word = 8'h10;
		16'h895D: out_word = 8'hF7;
		16'h895E: out_word = 8'hC9;
		16'h895F: out_word = 8'h46;
		16'h8960: out_word = 8'h23;
		16'h8961: out_word = 8'h7E;
		16'h8962: out_word = 8'hE5;
		16'h8963: out_word = 8'hC5;
		16'h8964: out_word = 8'hCD;
		16'h8965: out_word = 8'hA3;
		16'h8966: out_word = 8'h08;
		16'h8967: out_word = 8'hC1;
		16'h8968: out_word = 8'hE1;
		16'h8969: out_word = 8'h23;
		16'h896A: out_word = 8'h10;
		16'h896B: out_word = 8'hF5;
		16'h896C: out_word = 8'hC9;
		16'h896D: out_word = 8'hEF;
		16'h896E: out_word = 8'hAA;
		16'h896F: out_word = 8'h22;
		16'h8970: out_word = 8'h47;
		16'h8971: out_word = 8'h04;
		16'h8972: out_word = 8'hAF;
		16'h8973: out_word = 8'h37;
		16'h8974: out_word = 8'h1F;
		16'h8975: out_word = 8'h10;
		16'h8976: out_word = 8'hFD;
		16'h8977: out_word = 8'hA6;
		16'h8978: out_word = 8'hC9;
		16'h8979: out_word = 8'h06;
		16'h897A: out_word = 8'h1B;
		16'h897B: out_word = 8'h31;
		16'h897C: out_word = 8'h1B;
		16'h897D: out_word = 8'h4C;
		16'h897E: out_word = 8'h00;
		16'h897F: out_word = 8'h03;
		16'h8980: out_word = 8'h01;
		16'h8981: out_word = 8'h0A;
		16'h8982: out_word = 8'h02;
		16'h8983: out_word = 8'h1B;
		16'h8984: out_word = 8'h32;
		16'h8985: out_word = 8'hF3;
		16'h8986: out_word = 8'hC5;
		16'h8987: out_word = 8'h11;
		16'h8988: out_word = 8'h37;
		16'h8989: out_word = 8'h00;
		16'h898A: out_word = 8'h21;
		16'h898B: out_word = 8'h3C;
		16'h898C: out_word = 8'h00;
		16'h898D: out_word = 8'h19;
		16'h898E: out_word = 8'h10;
		16'h898F: out_word = 8'hFD;
		16'h8990: out_word = 8'h4D;
		16'h8991: out_word = 8'h44;
		16'h8992: out_word = 8'hEF;
		16'h8993: out_word = 8'h30;
		16'h8994: out_word = 8'h00;
		16'h8995: out_word = 8'hF3;
		16'h8996: out_word = 8'hD5;
		16'h8997: out_word = 8'hFD;
		16'h8998: out_word = 8'hE1;
		16'h8999: out_word = 8'hE5;
		16'h899A: out_word = 8'hDD;
		16'h899B: out_word = 8'hE1;
		16'h899C: out_word = 8'hFD;
		16'h899D: out_word = 8'h36;
		16'h899E: out_word = 8'h10;
		16'h899F: out_word = 8'hFF;
		16'h89A0: out_word = 8'h01;
		16'h89A1: out_word = 8'hC9;
		16'h89A2: out_word = 8'hFF;
		16'h89A3: out_word = 8'hDD;
		16'h89A4: out_word = 8'h09;
		16'h89A5: out_word = 8'hDD;
		16'h89A6: out_word = 8'h36;
		16'h89A7: out_word = 8'h03;
		16'h89A8: out_word = 8'h3C;
		16'h89A9: out_word = 8'hDD;
		16'h89AA: out_word = 8'h36;
		16'h89AB: out_word = 8'h01;
		16'h89AC: out_word = 8'hFF;
		16'h89AD: out_word = 8'hDD;
		16'h89AE: out_word = 8'h36;
		16'h89AF: out_word = 8'h04;
		16'h89B0: out_word = 8'h0F;
		16'h89B1: out_word = 8'hDD;
		16'h89B2: out_word = 8'h36;
		16'h89B3: out_word = 8'h05;
		16'h89B4: out_word = 8'h05;
		16'h89B5: out_word = 8'hDD;
		16'h89B6: out_word = 8'h36;
		16'h89B7: out_word = 8'h21;
		16'h89B8: out_word = 8'h00;
		16'h89B9: out_word = 8'hDD;
		16'h89BA: out_word = 8'h36;
		16'h89BB: out_word = 8'h0A;
		16'h89BC: out_word = 8'h00;
		16'h89BD: out_word = 8'hDD;
		16'h89BE: out_word = 8'h36;
		16'h89BF: out_word = 8'h0B;
		16'h89C0: out_word = 8'h00;
		16'h89C1: out_word = 8'hDD;
		16'h89C2: out_word = 8'h36;
		16'h89C3: out_word = 8'h16;
		16'h89C4: out_word = 8'hFF;
		16'h89C5: out_word = 8'hDD;
		16'h89C6: out_word = 8'h36;
		16'h89C7: out_word = 8'h17;
		16'h89C8: out_word = 8'h00;
		16'h89C9: out_word = 8'hDD;
		16'h89CA: out_word = 8'h36;
		16'h89CB: out_word = 8'h18;
		16'h89CC: out_word = 8'h00;
		16'h89CD: out_word = 8'hEF;
		16'h89CE: out_word = 8'hF1;
		16'h89CF: out_word = 8'h2B;
		16'h89D0: out_word = 8'hF3;
		16'h89D1: out_word = 8'hDD;
		16'h89D2: out_word = 8'h73;
		16'h89D3: out_word = 8'h06;
		16'h89D4: out_word = 8'hDD;
		16'h89D5: out_word = 8'h72;
		16'h89D6: out_word = 8'h07;
		16'h89D7: out_word = 8'hDD;
		16'h89D8: out_word = 8'h73;
		16'h89D9: out_word = 8'h0C;
		16'h89DA: out_word = 8'hDD;
		16'h89DB: out_word = 8'h72;
		16'h89DC: out_word = 8'h0D;
		16'h89DD: out_word = 8'hEB;
		16'h89DE: out_word = 8'h09;
		16'h89DF: out_word = 8'hDD;
		16'h89E0: out_word = 8'h75;
		16'h89E1: out_word = 8'h08;
		16'h89E2: out_word = 8'hDD;
		16'h89E3: out_word = 8'h74;
		16'h89E4: out_word = 8'h09;
		16'h89E5: out_word = 8'hC1;
		16'h89E6: out_word = 8'hC5;
		16'h89E7: out_word = 8'h05;
		16'h89E8: out_word = 8'h48;
		16'h89E9: out_word = 8'h06;
		16'h89EA: out_word = 8'h00;
		16'h89EB: out_word = 8'hCB;
		16'h89EC: out_word = 8'h21;
		16'h89ED: out_word = 8'hFD;
		16'h89EE: out_word = 8'hE5;
		16'h89EF: out_word = 8'hE1;
		16'h89F0: out_word = 8'h09;
		16'h89F1: out_word = 8'hDD;
		16'h89F2: out_word = 8'hE5;
		16'h89F3: out_word = 8'hC1;
		16'h89F4: out_word = 8'h71;
		16'h89F5: out_word = 8'h23;
		16'h89F6: out_word = 8'h70;
		16'h89F7: out_word = 8'hB7;
		16'h89F8: out_word = 8'hFD;
		16'h89F9: out_word = 8'hCB;
		16'h89FA: out_word = 8'h10;
		16'h89FB: out_word = 8'h16;
		16'h89FC: out_word = 8'hC1;
		16'h89FD: out_word = 8'h05;
		16'h89FE: out_word = 8'hC5;
		16'h89FF: out_word = 8'hDD;
		16'h8A00: out_word = 8'h70;
		16'h8A01: out_word = 8'h02;
		16'h8A02: out_word = 8'h20;
		16'h8A03: out_word = 8'h9C;
		16'h8A04: out_word = 8'hC1;
		16'h8A05: out_word = 8'hFD;
		16'h8A06: out_word = 8'h36;
		16'h8A07: out_word = 8'h27;
		16'h8A08: out_word = 8'h1A;
		16'h8A09: out_word = 8'hFD;
		16'h8A0A: out_word = 8'h36;
		16'h8A0B: out_word = 8'h28;
		16'h8A0C: out_word = 8'h0B;
		16'h8A0D: out_word = 8'hFD;
		16'h8A0E: out_word = 8'hE5;
		16'h8A0F: out_word = 8'hE1;
		16'h8A10: out_word = 8'h01;
		16'h8A11: out_word = 8'h2B;
		16'h8A12: out_word = 8'h00;
		16'h8A13: out_word = 8'h09;
		16'h8A14: out_word = 8'hEB;
		16'h8A15: out_word = 8'h21;
		16'h8A16: out_word = 8'h31;
		16'h8A17: out_word = 8'h0A;
		16'h8A18: out_word = 8'h01;
		16'h8A19: out_word = 8'h0D;
		16'h8A1A: out_word = 8'h00;
		16'h8A1B: out_word = 8'hED;
		16'h8A1C: out_word = 8'hB0;
		16'h8A1D: out_word = 8'h16;
		16'h8A1E: out_word = 8'h07;
		16'h8A1F: out_word = 8'h1E;
		16'h8A20: out_word = 8'hF8;
		16'h8A21: out_word = 8'hCD;
		16'h8A22: out_word = 8'h7C;
		16'h8A23: out_word = 8'h0E;
		16'h8A24: out_word = 8'h16;
		16'h8A25: out_word = 8'h0B;
		16'h8A26: out_word = 8'h1E;
		16'h8A27: out_word = 8'hFF;
		16'h8A28: out_word = 8'hCD;
		16'h8A29: out_word = 8'h7C;
		16'h8A2A: out_word = 8'h0E;
		16'h8A2B: out_word = 8'h14;
		16'h8A2C: out_word = 8'hCD;
		16'h8A2D: out_word = 8'h7C;
		16'h8A2E: out_word = 8'h0E;
		16'h8A2F: out_word = 8'h18;
		16'h8A30: out_word = 8'h4C;
		16'h8A31: out_word = 8'hEF;
		16'h8A32: out_word = 8'hA4;
		16'h8A33: out_word = 8'h01;
		16'h8A34: out_word = 8'h05;
		16'h8A35: out_word = 8'h34;
		16'h8A36: out_word = 8'hDF;
		16'h8A37: out_word = 8'h75;
		16'h8A38: out_word = 8'hF4;
		16'h8A39: out_word = 8'h38;
		16'h8A3A: out_word = 8'h75;
		16'h8A3B: out_word = 8'h05;
		16'h8A3C: out_word = 8'h38;
		16'h8A3D: out_word = 8'hC9;
		16'h8A3E: out_word = 8'h3E;
		16'h8A3F: out_word = 8'h7F;
		16'h8A40: out_word = 8'hDB;
		16'h8A41: out_word = 8'hFE;
		16'h8A42: out_word = 8'h1F;
		16'h8A43: out_word = 8'hD8;
		16'h8A44: out_word = 8'h3E;
		16'h8A45: out_word = 8'hFE;
		16'h8A46: out_word = 8'hDB;
		16'h8A47: out_word = 8'hFE;
		16'h8A48: out_word = 8'h1F;
		16'h8A49: out_word = 8'hC9;
		16'h8A4A: out_word = 8'h01;
		16'h8A4B: out_word = 8'h11;
		16'h8A4C: out_word = 8'h00;
		16'h8A4D: out_word = 8'h18;
		16'h8A4E: out_word = 8'h03;
		16'h8A4F: out_word = 8'h01;
		16'h8A50: out_word = 8'h00;
		16'h8A51: out_word = 8'h00;
		16'h8A52: out_word = 8'hFD;
		16'h8A53: out_word = 8'hE5;
		16'h8A54: out_word = 8'hE1;
		16'h8A55: out_word = 8'h09;
		16'h8A56: out_word = 8'hFD;
		16'h8A57: out_word = 8'h75;
		16'h8A58: out_word = 8'h23;
		16'h8A59: out_word = 8'hFD;
		16'h8A5A: out_word = 8'h74;
		16'h8A5B: out_word = 8'h24;
		16'h8A5C: out_word = 8'hFD;
		16'h8A5D: out_word = 8'h7E;
		16'h8A5E: out_word = 8'h10;
		16'h8A5F: out_word = 8'hFD;
		16'h8A60: out_word = 8'h77;
		16'h8A61: out_word = 8'h22;
		16'h8A62: out_word = 8'hFD;
		16'h8A63: out_word = 8'h36;
		16'h8A64: out_word = 8'h21;
		16'h8A65: out_word = 8'h01;
		16'h8A66: out_word = 8'hC9;
		16'h8A67: out_word = 8'h5E;
		16'h8A68: out_word = 8'h23;
		16'h8A69: out_word = 8'h56;
		16'h8A6A: out_word = 8'hD5;
		16'h8A6B: out_word = 8'hDD;
		16'h8A6C: out_word = 8'hE1;
		16'h8A6D: out_word = 8'hC9;
		16'h8A6E: out_word = 8'hFD;
		16'h8A6F: out_word = 8'h6E;
		16'h8A70: out_word = 8'h23;
		16'h8A71: out_word = 8'hFD;
		16'h8A72: out_word = 8'h66;
		16'h8A73: out_word = 8'h24;
		16'h8A74: out_word = 8'h23;
		16'h8A75: out_word = 8'h23;
		16'h8A76: out_word = 8'hFD;
		16'h8A77: out_word = 8'h75;
		16'h8A78: out_word = 8'h23;
		16'h8A79: out_word = 8'hFD;
		16'h8A7A: out_word = 8'h74;
		16'h8A7B: out_word = 8'h24;
		16'h8A7C: out_word = 8'hC9;
		16'h8A7D: out_word = 8'hCD;
		16'h8A7E: out_word = 8'h4F;
		16'h8A7F: out_word = 8'h0A;
		16'h8A80: out_word = 8'hFD;
		16'h8A81: out_word = 8'hCB;
		16'h8A82: out_word = 8'h22;
		16'h8A83: out_word = 8'h1E;
		16'h8A84: out_word = 8'h38;
		16'h8A85: out_word = 8'h06;
		16'h8A86: out_word = 8'hCD;
		16'h8A87: out_word = 8'h67;
		16'h8A88: out_word = 8'h0A;
		16'h8A89: out_word = 8'hCD;
		16'h8A8A: out_word = 8'h5C;
		16'h8A8B: out_word = 8'h0B;
		16'h8A8C: out_word = 8'hFD;
		16'h8A8D: out_word = 8'hCB;
		16'h8A8E: out_word = 8'h21;
		16'h8A8F: out_word = 8'h26;
		16'h8A90: out_word = 8'h38;
		16'h8A91: out_word = 8'h05;
		16'h8A92: out_word = 8'hCD;
		16'h8A93: out_word = 8'h6E;
		16'h8A94: out_word = 8'h0A;
		16'h8A95: out_word = 8'h18;
		16'h8A96: out_word = 8'hE9;
		16'h8A97: out_word = 8'hCD;
		16'h8A98: out_word = 8'h91;
		16'h8A99: out_word = 8'h0F;
		16'h8A9A: out_word = 8'hD5;
		16'h8A9B: out_word = 8'hCD;
		16'h8A9C: out_word = 8'h42;
		16'h8A9D: out_word = 8'h0F;
		16'h8A9E: out_word = 8'hD1;
		16'h8A9F: out_word = 8'hFD;
		16'h8AA0: out_word = 8'h7E;
		16'h8AA1: out_word = 8'h10;
		16'h8AA2: out_word = 8'hFE;
		16'h8AA3: out_word = 8'hFF;
		16'h8AA4: out_word = 8'h20;
		16'h8AA5: out_word = 8'h05;
		16'h8AA6: out_word = 8'hCD;
		16'h8AA7: out_word = 8'h93;
		16'h8AA8: out_word = 8'h0E;
		16'h8AA9: out_word = 8'hFB;
		16'h8AAA: out_word = 8'hC9;
		16'h8AAB: out_word = 8'h1B;
		16'h8AAC: out_word = 8'hCD;
		16'h8AAD: out_word = 8'h76;
		16'h8AAE: out_word = 8'h0F;
		16'h8AAF: out_word = 8'hCD;
		16'h8AB0: out_word = 8'hC1;
		16'h8AB1: out_word = 8'h0F;
		16'h8AB2: out_word = 8'hCD;
		16'h8AB3: out_word = 8'h91;
		16'h8AB4: out_word = 8'h0F;
		16'h8AB5: out_word = 8'h18;
		16'h8AB6: out_word = 8'hE8;
		16'h8AB7: out_word = 8'h48;
		16'h8AB8: out_word = 8'h5A;
		16'h8AB9: out_word = 8'h59;
		16'h8ABA: out_word = 8'h58;
		16'h8ABB: out_word = 8'h57;
		16'h8ABC: out_word = 8'h55;
		16'h8ABD: out_word = 8'h56;
		16'h8ABE: out_word = 8'h4D;
		16'h8ABF: out_word = 8'h54;
		16'h8AC0: out_word = 8'h29;
		16'h8AC1: out_word = 8'h28;
		16'h8AC2: out_word = 8'h4E;
		16'h8AC3: out_word = 8'h4F;
		16'h8AC4: out_word = 8'h21;
		16'h8AC5: out_word = 8'hCD;
		16'h8AC6: out_word = 8'hE3;
		16'h8AC7: out_word = 8'h0E;
		16'h8AC8: out_word = 8'hD8;
		16'h8AC9: out_word = 8'hDD;
		16'h8ACA: out_word = 8'h34;
		16'h8ACB: out_word = 8'h06;
		16'h8ACC: out_word = 8'hC0;
		16'h8ACD: out_word = 8'hDD;
		16'h8ACE: out_word = 8'h34;
		16'h8ACF: out_word = 8'h07;
		16'h8AD0: out_word = 8'hC9;
		16'h8AD1: out_word = 8'hE5;
		16'h8AD2: out_word = 8'h0E;
		16'h8AD3: out_word = 8'h00;
		16'h8AD4: out_word = 8'hCD;
		16'h8AD5: out_word = 8'hC5;
		16'h8AD6: out_word = 8'h0A;
		16'h8AD7: out_word = 8'h38;
		16'h8AD8: out_word = 8'h08;
		16'h8AD9: out_word = 8'hFE;
		16'h8ADA: out_word = 8'h26;
		16'h8ADB: out_word = 8'h20;
		16'h8ADC: out_word = 8'h0F;
		16'h8ADD: out_word = 8'h3E;
		16'h8ADE: out_word = 8'h80;
		16'h8ADF: out_word = 8'hE1;
		16'h8AE0: out_word = 8'hC9;
		16'h8AE1: out_word = 8'hFD;
		16'h8AE2: out_word = 8'h7E;
		16'h8AE3: out_word = 8'h21;
		16'h8AE4: out_word = 8'hFD;
		16'h8AE5: out_word = 8'hB6;
		16'h8AE6: out_word = 8'h10;
		16'h8AE7: out_word = 8'hFD;
		16'h8AE8: out_word = 8'h77;
		16'h8AE9: out_word = 8'h10;
		16'h8AEA: out_word = 8'h18;
		16'h8AEB: out_word = 8'hF3;
		16'h8AEC: out_word = 8'hFE;
		16'h8AED: out_word = 8'h23;
		16'h8AEE: out_word = 8'h20;
		16'h8AEF: out_word = 8'h03;
		16'h8AF0: out_word = 8'h0C;
		16'h8AF1: out_word = 8'h18;
		16'h8AF2: out_word = 8'hE1;
		16'h8AF3: out_word = 8'hFE;
		16'h8AF4: out_word = 8'h24;
		16'h8AF5: out_word = 8'h20;
		16'h8AF6: out_word = 8'h03;
		16'h8AF7: out_word = 8'h0D;
		16'h8AF8: out_word = 8'h18;
		16'h8AF9: out_word = 8'hDA;
		16'h8AFA: out_word = 8'hCB;
		16'h8AFB: out_word = 8'h6F;
		16'h8AFC: out_word = 8'h20;
		16'h8AFD: out_word = 8'h06;
		16'h8AFE: out_word = 8'hF5;
		16'h8AFF: out_word = 8'h3E;
		16'h8B00: out_word = 8'h0C;
		16'h8B01: out_word = 8'h81;
		16'h8B02: out_word = 8'h4F;
		16'h8B03: out_word = 8'hF1;
		16'h8B04: out_word = 8'hE6;
		16'h8B05: out_word = 8'hDF;
		16'h8B06: out_word = 8'hD6;
		16'h8B07: out_word = 8'h41;
		16'h8B08: out_word = 8'hDA;
		16'h8B09: out_word = 8'h22;
		16'h8B0A: out_word = 8'h0F;
		16'h8B0B: out_word = 8'hFE;
		16'h8B0C: out_word = 8'h07;
		16'h8B0D: out_word = 8'hD2;
		16'h8B0E: out_word = 8'h22;
		16'h8B0F: out_word = 8'h0F;
		16'h8B10: out_word = 8'hC5;
		16'h8B11: out_word = 8'h06;
		16'h8B12: out_word = 8'h00;
		16'h8B13: out_word = 8'h4F;
		16'h8B14: out_word = 8'h21;
		16'h8B15: out_word = 8'hF9;
		16'h8B16: out_word = 8'h0D;
		16'h8B17: out_word = 8'h09;
		16'h8B18: out_word = 8'h7E;
		16'h8B19: out_word = 8'hC1;
		16'h8B1A: out_word = 8'h81;
		16'h8B1B: out_word = 8'hE1;
		16'h8B1C: out_word = 8'hC9;
		16'h8B1D: out_word = 8'hE5;
		16'h8B1E: out_word = 8'hD5;
		16'h8B1F: out_word = 8'hDD;
		16'h8B20: out_word = 8'h6E;
		16'h8B21: out_word = 8'h06;
		16'h8B22: out_word = 8'hDD;
		16'h8B23: out_word = 8'h66;
		16'h8B24: out_word = 8'h07;
		16'h8B25: out_word = 8'h11;
		16'h8B26: out_word = 8'h00;
		16'h8B27: out_word = 8'h00;
		16'h8B28: out_word = 8'h7E;
		16'h8B29: out_word = 8'hFE;
		16'h8B2A: out_word = 8'h30;
		16'h8B2B: out_word = 8'h38;
		16'h8B2C: out_word = 8'h18;
		16'h8B2D: out_word = 8'hFE;
		16'h8B2E: out_word = 8'h3A;
		16'h8B2F: out_word = 8'h30;
		16'h8B30: out_word = 8'h14;
		16'h8B31: out_word = 8'h23;
		16'h8B32: out_word = 8'hE5;
		16'h8B33: out_word = 8'hCD;
		16'h8B34: out_word = 8'h50;
		16'h8B35: out_word = 8'h0B;
		16'h8B36: out_word = 8'hD6;
		16'h8B37: out_word = 8'h30;
		16'h8B38: out_word = 8'h26;
		16'h8B39: out_word = 8'h00;
		16'h8B3A: out_word = 8'h6F;
		16'h8B3B: out_word = 8'h19;
		16'h8B3C: out_word = 8'h38;
		16'h8B3D: out_word = 8'h04;
		16'h8B3E: out_word = 8'hEB;
		16'h8B3F: out_word = 8'hE1;
		16'h8B40: out_word = 8'h18;
		16'h8B41: out_word = 8'hE6;
		16'h8B42: out_word = 8'hC3;
		16'h8B43: out_word = 8'h1A;
		16'h8B44: out_word = 8'h0F;
		16'h8B45: out_word = 8'hDD;
		16'h8B46: out_word = 8'h75;
		16'h8B47: out_word = 8'h06;
		16'h8B48: out_word = 8'hDD;
		16'h8B49: out_word = 8'h74;
		16'h8B4A: out_word = 8'h07;
		16'h8B4B: out_word = 8'hD5;
		16'h8B4C: out_word = 8'hC1;
		16'h8B4D: out_word = 8'hD1;
		16'h8B4E: out_word = 8'hE1;
		16'h8B4F: out_word = 8'hC9;
		16'h8B50: out_word = 8'h21;
		16'h8B51: out_word = 8'h00;
		16'h8B52: out_word = 8'h00;
		16'h8B53: out_word = 8'h06;
		16'h8B54: out_word = 8'h0A;
		16'h8B55: out_word = 8'h19;
		16'h8B56: out_word = 8'h38;
		16'h8B57: out_word = 8'hEA;
		16'h8B58: out_word = 8'h10;
		16'h8B59: out_word = 8'hFB;
		16'h8B5A: out_word = 8'hEB;
		16'h8B5B: out_word = 8'hC9;
		16'h8B5C: out_word = 8'hCD;
		16'h8B5D: out_word = 8'h3E;
		16'h8B5E: out_word = 8'h0A;
		16'h8B5F: out_word = 8'h38;
		16'h8B60: out_word = 8'h08;
		16'h8B61: out_word = 8'hCD;
		16'h8B62: out_word = 8'h93;
		16'h8B63: out_word = 8'h0E;
		16'h8B64: out_word = 8'hFB;
		16'h8B65: out_word = 8'hCD;
		16'h8B66: out_word = 8'hAC;
		16'h8B67: out_word = 8'h05;
		16'h8B68: out_word = 8'h14;
		16'h8B69: out_word = 8'hCD;
		16'h8B6A: out_word = 8'hC5;
		16'h8B6B: out_word = 8'h0A;
		16'h8B6C: out_word = 8'hDA;
		16'h8B6D: out_word = 8'hA2;
		16'h8B6E: out_word = 8'h0D;
		16'h8B6F: out_word = 8'hCD;
		16'h8B70: out_word = 8'hF0;
		16'h8B71: out_word = 8'h0D;
		16'h8B72: out_word = 8'h06;
		16'h8B73: out_word = 8'h00;
		16'h8B74: out_word = 8'hCB;
		16'h8B75: out_word = 8'h21;
		16'h8B76: out_word = 8'h21;
		16'h8B77: out_word = 8'hCA;
		16'h8B78: out_word = 8'h0D;
		16'h8B79: out_word = 8'h09;
		16'h8B7A: out_word = 8'h5E;
		16'h8B7B: out_word = 8'h23;
		16'h8B7C: out_word = 8'h56;
		16'h8B7D: out_word = 8'hEB;
		16'h8B7E: out_word = 8'hCD;
		16'h8B7F: out_word = 8'h84;
		16'h8B80: out_word = 8'h0B;
		16'h8B81: out_word = 8'h18;
		16'h8B82: out_word = 8'hD9;
		16'h8B83: out_word = 8'hC9;
		16'h8B84: out_word = 8'hE9;
		16'h8B85: out_word = 8'hCD;
		16'h8B86: out_word = 8'hC5;
		16'h8B87: out_word = 8'h0A;
		16'h8B88: out_word = 8'hDA;
		16'h8B89: out_word = 8'hA1;
		16'h8B8A: out_word = 8'h0D;
		16'h8B8B: out_word = 8'hFE;
		16'h8B8C: out_word = 8'h21;
		16'h8B8D: out_word = 8'hC8;
		16'h8B8E: out_word = 8'h18;
		16'h8B8F: out_word = 8'hF5;
		16'h8B90: out_word = 8'hCD;
		16'h8B91: out_word = 8'h1D;
		16'h8B92: out_word = 8'h0B;
		16'h8B93: out_word = 8'h79;
		16'h8B94: out_word = 8'hFE;
		16'h8B95: out_word = 8'h09;
		16'h8B96: out_word = 8'hD2;
		16'h8B97: out_word = 8'h12;
		16'h8B98: out_word = 8'h0F;
		16'h8B99: out_word = 8'hCB;
		16'h8B9A: out_word = 8'h27;
		16'h8B9B: out_word = 8'hCB;
		16'h8B9C: out_word = 8'h27;
		16'h8B9D: out_word = 8'h47;
		16'h8B9E: out_word = 8'hCB;
		16'h8B9F: out_word = 8'h27;
		16'h8BA0: out_word = 8'h80;
		16'h8BA1: out_word = 8'hDD;
		16'h8BA2: out_word = 8'h77;
		16'h8BA3: out_word = 8'h03;
		16'h8BA4: out_word = 8'hC9;
		16'h8BA5: out_word = 8'hC9;
		16'h8BA6: out_word = 8'hDD;
		16'h8BA7: out_word = 8'h7E;
		16'h8BA8: out_word = 8'h0B;
		16'h8BA9: out_word = 8'h3C;
		16'h8BAA: out_word = 8'hFE;
		16'h8BAB: out_word = 8'h05;
		16'h8BAC: out_word = 8'hCA;
		16'h8BAD: out_word = 8'h2A;
		16'h8BAE: out_word = 8'h0F;
		16'h8BAF: out_word = 8'hDD;
		16'h8BB0: out_word = 8'h77;
		16'h8BB1: out_word = 8'h0B;
		16'h8BB2: out_word = 8'h11;
		16'h8BB3: out_word = 8'h0C;
		16'h8BB4: out_word = 8'h00;
		16'h8BB5: out_word = 8'hCD;
		16'h8BB6: out_word = 8'h27;
		16'h8BB7: out_word = 8'h0C;
		16'h8BB8: out_word = 8'hDD;
		16'h8BB9: out_word = 8'h7E;
		16'h8BBA: out_word = 8'h06;
		16'h8BBB: out_word = 8'h77;
		16'h8BBC: out_word = 8'h23;
		16'h8BBD: out_word = 8'hDD;
		16'h8BBE: out_word = 8'h7E;
		16'h8BBF: out_word = 8'h07;
		16'h8BC0: out_word = 8'h77;
		16'h8BC1: out_word = 8'hC9;
		16'h8BC2: out_word = 8'hDD;
		16'h8BC3: out_word = 8'h7E;
		16'h8BC4: out_word = 8'h16;
		16'h8BC5: out_word = 8'h11;
		16'h8BC6: out_word = 8'h17;
		16'h8BC7: out_word = 8'h00;
		16'h8BC8: out_word = 8'hB7;
		16'h8BC9: out_word = 8'hFA;
		16'h8BCA: out_word = 8'hF0;
		16'h8BCB: out_word = 8'h0B;
		16'h8BCC: out_word = 8'hCD;
		16'h8BCD: out_word = 8'h27;
		16'h8BCE: out_word = 8'h0C;
		16'h8BCF: out_word = 8'hDD;
		16'h8BD0: out_word = 8'h7E;
		16'h8BD1: out_word = 8'h06;
		16'h8BD2: out_word = 8'hBE;
		16'h8BD3: out_word = 8'h20;
		16'h8BD4: out_word = 8'h1B;
		16'h8BD5: out_word = 8'h23;
		16'h8BD6: out_word = 8'hDD;
		16'h8BD7: out_word = 8'h7E;
		16'h8BD8: out_word = 8'h07;
		16'h8BD9: out_word = 8'hBE;
		16'h8BDA: out_word = 8'h20;
		16'h8BDB: out_word = 8'h14;
		16'h8BDC: out_word = 8'hDD;
		16'h8BDD: out_word = 8'h35;
		16'h8BDE: out_word = 8'h16;
		16'h8BDF: out_word = 8'hDD;
		16'h8BE0: out_word = 8'h7E;
		16'h8BE1: out_word = 8'h16;
		16'h8BE2: out_word = 8'hB7;
		16'h8BE3: out_word = 8'hF0;
		16'h8BE4: out_word = 8'hDD;
		16'h8BE5: out_word = 8'hCB;
		16'h8BE6: out_word = 8'h0A;
		16'h8BE7: out_word = 8'h46;
		16'h8BE8: out_word = 8'hC8;
		16'h8BE9: out_word = 8'hDD;
		16'h8BEA: out_word = 8'h36;
		16'h8BEB: out_word = 8'h16;
		16'h8BEC: out_word = 8'h00;
		16'h8BED: out_word = 8'hAF;
		16'h8BEE: out_word = 8'h18;
		16'h8BEF: out_word = 8'h1B;
		16'h8BF0: out_word = 8'hDD;
		16'h8BF1: out_word = 8'h7E;
		16'h8BF2: out_word = 8'h16;
		16'h8BF3: out_word = 8'h3C;
		16'h8BF4: out_word = 8'hFE;
		16'h8BF5: out_word = 8'h05;
		16'h8BF6: out_word = 8'hCA;
		16'h8BF7: out_word = 8'h2A;
		16'h8BF8: out_word = 8'h0F;
		16'h8BF9: out_word = 8'hDD;
		16'h8BFA: out_word = 8'h77;
		16'h8BFB: out_word = 8'h16;
		16'h8BFC: out_word = 8'hCD;
		16'h8BFD: out_word = 8'h27;
		16'h8BFE: out_word = 8'h0C;
		16'h8BFF: out_word = 8'hDD;
		16'h8C00: out_word = 8'h7E;
		16'h8C01: out_word = 8'h06;
		16'h8C02: out_word = 8'h77;
		16'h8C03: out_word = 8'h23;
		16'h8C04: out_word = 8'hDD;
		16'h8C05: out_word = 8'h7E;
		16'h8C06: out_word = 8'h07;
		16'h8C07: out_word = 8'h77;
		16'h8C08: out_word = 8'hDD;
		16'h8C09: out_word = 8'h7E;
		16'h8C0A: out_word = 8'h0B;
		16'h8C0B: out_word = 8'h11;
		16'h8C0C: out_word = 8'h0C;
		16'h8C0D: out_word = 8'h00;
		16'h8C0E: out_word = 8'hCD;
		16'h8C0F: out_word = 8'h27;
		16'h8C10: out_word = 8'h0C;
		16'h8C11: out_word = 8'h7E;
		16'h8C12: out_word = 8'hDD;
		16'h8C13: out_word = 8'h77;
		16'h8C14: out_word = 8'h06;
		16'h8C15: out_word = 8'h23;
		16'h8C16: out_word = 8'h7E;
		16'h8C17: out_word = 8'hDD;
		16'h8C18: out_word = 8'h77;
		16'h8C19: out_word = 8'h07;
		16'h8C1A: out_word = 8'hDD;
		16'h8C1B: out_word = 8'h35;
		16'h8C1C: out_word = 8'h0B;
		16'h8C1D: out_word = 8'hF0;
		16'h8C1E: out_word = 8'hDD;
		16'h8C1F: out_word = 8'h36;
		16'h8C20: out_word = 8'h0B;
		16'h8C21: out_word = 8'h00;
		16'h8C22: out_word = 8'hDD;
		16'h8C23: out_word = 8'hCB;
		16'h8C24: out_word = 8'h0A;
		16'h8C25: out_word = 8'hC6;
		16'h8C26: out_word = 8'hC9;
		16'h8C27: out_word = 8'hDD;
		16'h8C28: out_word = 8'hE5;
		16'h8C29: out_word = 8'hE1;
		16'h8C2A: out_word = 8'h19;
		16'h8C2B: out_word = 8'h06;
		16'h8C2C: out_word = 8'h00;
		16'h8C2D: out_word = 8'h4F;
		16'h8C2E: out_word = 8'hCB;
		16'h8C2F: out_word = 8'h21;
		16'h8C30: out_word = 8'h09;
		16'h8C31: out_word = 8'hC9;
		16'h8C32: out_word = 8'hCD;
		16'h8C33: out_word = 8'h1D;
		16'h8C34: out_word = 8'h0B;
		16'h8C35: out_word = 8'h78;
		16'h8C36: out_word = 8'hB7;
		16'h8C37: out_word = 8'hC2;
		16'h8C38: out_word = 8'h12;
		16'h8C39: out_word = 8'h0F;
		16'h8C3A: out_word = 8'h79;
		16'h8C3B: out_word = 8'hFE;
		16'h8C3C: out_word = 8'h3C;
		16'h8C3D: out_word = 8'hDA;
		16'h8C3E: out_word = 8'h12;
		16'h8C3F: out_word = 8'h0F;
		16'h8C40: out_word = 8'hFE;
		16'h8C41: out_word = 8'hF1;
		16'h8C42: out_word = 8'hD2;
		16'h8C43: out_word = 8'h12;
		16'h8C44: out_word = 8'h0F;
		16'h8C45: out_word = 8'hDD;
		16'h8C46: out_word = 8'h7E;
		16'h8C47: out_word = 8'h02;
		16'h8C48: out_word = 8'hB7;
		16'h8C49: out_word = 8'hC0;
		16'h8C4A: out_word = 8'h06;
		16'h8C4B: out_word = 8'h00;
		16'h8C4C: out_word = 8'hC5;
		16'h8C4D: out_word = 8'hE1;
		16'h8C4E: out_word = 8'h29;
		16'h8C4F: out_word = 8'h29;
		16'h8C50: out_word = 8'hE5;
		16'h8C51: out_word = 8'hC1;
		16'h8C52: out_word = 8'hFD;
		16'h8C53: out_word = 8'hE5;
		16'h8C54: out_word = 8'hEF;
		16'h8C55: out_word = 8'h2B;
		16'h8C56: out_word = 8'h2D;
		16'h8C57: out_word = 8'hF3;
		16'h8C58: out_word = 8'hFD;
		16'h8C59: out_word = 8'hE1;
		16'h8C5A: out_word = 8'hFD;
		16'h8C5B: out_word = 8'hE5;
		16'h8C5C: out_word = 8'hFD;
		16'h8C5D: out_word = 8'hE5;
		16'h8C5E: out_word = 8'hE1;
		16'h8C5F: out_word = 8'h01;
		16'h8C60: out_word = 8'h2B;
		16'h8C61: out_word = 8'h00;
		16'h8C62: out_word = 8'h09;
		16'h8C63: out_word = 8'hFD;
		16'h8C64: out_word = 8'h21;
		16'h8C65: out_word = 8'h3A;
		16'h8C66: out_word = 8'h5C;
		16'h8C67: out_word = 8'hE5;
		16'h8C68: out_word = 8'h21;
		16'h8C69: out_word = 8'h76;
		16'h8C6A: out_word = 8'h0C;
		16'h8C6B: out_word = 8'h22;
		16'h8C6C: out_word = 8'h5A;
		16'h8C6D: out_word = 8'h5B;
		16'h8C6E: out_word = 8'h21;
		16'h8C6F: out_word = 8'h14;
		16'h8C70: out_word = 8'h5B;
		16'h8C71: out_word = 8'hE3;
		16'h8C72: out_word = 8'hE5;
		16'h8C73: out_word = 8'hC3;
		16'h8C74: out_word = 8'h00;
		16'h8C75: out_word = 8'h5B;
		16'h8C76: out_word = 8'hF3;
		16'h8C77: out_word = 8'hEF;
		16'h8C78: out_word = 8'hA2;
		16'h8C79: out_word = 8'h2D;
		16'h8C7A: out_word = 8'hF3;
		16'h8C7B: out_word = 8'hFD;
		16'h8C7C: out_word = 8'hE1;
		16'h8C7D: out_word = 8'hFD;
		16'h8C7E: out_word = 8'h71;
		16'h8C7F: out_word = 8'h27;
		16'h8C80: out_word = 8'hFD;
		16'h8C81: out_word = 8'h70;
		16'h8C82: out_word = 8'h28;
		16'h8C83: out_word = 8'hC9;
		16'h8C84: out_word = 8'hCD;
		16'h8C85: out_word = 8'h1D;
		16'h8C86: out_word = 8'h0B;
		16'h8C87: out_word = 8'h79;
		16'h8C88: out_word = 8'hFE;
		16'h8C89: out_word = 8'h40;
		16'h8C8A: out_word = 8'hD2;
		16'h8C8B: out_word = 8'h12;
		16'h8C8C: out_word = 8'h0F;
		16'h8C8D: out_word = 8'h2F;
		16'h8C8E: out_word = 8'h5F;
		16'h8C8F: out_word = 8'h16;
		16'h8C90: out_word = 8'h07;
		16'h8C91: out_word = 8'hCD;
		16'h8C92: out_word = 8'h7C;
		16'h8C93: out_word = 8'h0E;
		16'h8C94: out_word = 8'hC9;
		16'h8C95: out_word = 8'hCD;
		16'h8C96: out_word = 8'h1D;
		16'h8C97: out_word = 8'h0B;
		16'h8C98: out_word = 8'h79;
		16'h8C99: out_word = 8'hFE;
		16'h8C9A: out_word = 8'h10;
		16'h8C9B: out_word = 8'hD2;
		16'h8C9C: out_word = 8'h12;
		16'h8C9D: out_word = 8'h0F;
		16'h8C9E: out_word = 8'hDD;
		16'h8C9F: out_word = 8'h77;
		16'h8CA0: out_word = 8'h04;
		16'h8CA1: out_word = 8'hDD;
		16'h8CA2: out_word = 8'h5E;
		16'h8CA3: out_word = 8'h02;
		16'h8CA4: out_word = 8'h3E;
		16'h8CA5: out_word = 8'h08;
		16'h8CA6: out_word = 8'h83;
		16'h8CA7: out_word = 8'h57;
		16'h8CA8: out_word = 8'h59;
		16'h8CA9: out_word = 8'hCD;
		16'h8CAA: out_word = 8'h7C;
		16'h8CAB: out_word = 8'h0E;
		16'h8CAC: out_word = 8'hC9;
		16'h8CAD: out_word = 8'hDD;
		16'h8CAE: out_word = 8'h5E;
		16'h8CAF: out_word = 8'h02;
		16'h8CB0: out_word = 8'h3E;
		16'h8CB1: out_word = 8'h08;
		16'h8CB2: out_word = 8'h83;
		16'h8CB3: out_word = 8'h57;
		16'h8CB4: out_word = 8'h1E;
		16'h8CB5: out_word = 8'h1F;
		16'h8CB6: out_word = 8'hDD;
		16'h8CB7: out_word = 8'h73;
		16'h8CB8: out_word = 8'h04;
		16'h8CB9: out_word = 8'hC9;
		16'h8CBA: out_word = 8'hCD;
		16'h8CBB: out_word = 8'h1D;
		16'h8CBC: out_word = 8'h0B;
		16'h8CBD: out_word = 8'h79;
		16'h8CBE: out_word = 8'hFE;
		16'h8CBF: out_word = 8'h08;
		16'h8CC0: out_word = 8'hD2;
		16'h8CC1: out_word = 8'h12;
		16'h8CC2: out_word = 8'h0F;
		16'h8CC3: out_word = 8'h06;
		16'h8CC4: out_word = 8'h00;
		16'h8CC5: out_word = 8'h21;
		16'h8CC6: out_word = 8'hE8;
		16'h8CC7: out_word = 8'h0D;
		16'h8CC8: out_word = 8'h09;
		16'h8CC9: out_word = 8'h7E;
		16'h8CCA: out_word = 8'hFD;
		16'h8CCB: out_word = 8'h77;
		16'h8CCC: out_word = 8'h29;
		16'h8CCD: out_word = 8'hC9;
		16'h8CCE: out_word = 8'hCD;
		16'h8CCF: out_word = 8'h1D;
		16'h8CD0: out_word = 8'h0B;
		16'h8CD1: out_word = 8'h16;
		16'h8CD2: out_word = 8'h0B;
		16'h8CD3: out_word = 8'h59;
		16'h8CD4: out_word = 8'hCD;
		16'h8CD5: out_word = 8'h7C;
		16'h8CD6: out_word = 8'h0E;
		16'h8CD7: out_word = 8'h14;
		16'h8CD8: out_word = 8'h58;
		16'h8CD9: out_word = 8'hCD;
		16'h8CDA: out_word = 8'h7C;
		16'h8CDB: out_word = 8'h0E;
		16'h8CDC: out_word = 8'hC9;
		16'h8CDD: out_word = 8'hCD;
		16'h8CDE: out_word = 8'h1D;
		16'h8CDF: out_word = 8'h0B;
		16'h8CE0: out_word = 8'h79;
		16'h8CE1: out_word = 8'h3D;
		16'h8CE2: out_word = 8'hFA;
		16'h8CE3: out_word = 8'h12;
		16'h8CE4: out_word = 8'h0F;
		16'h8CE5: out_word = 8'hFE;
		16'h8CE6: out_word = 8'h10;
		16'h8CE7: out_word = 8'hD2;
		16'h8CE8: out_word = 8'h12;
		16'h8CE9: out_word = 8'h0F;
		16'h8CEA: out_word = 8'hDD;
		16'h8CEB: out_word = 8'h77;
		16'h8CEC: out_word = 8'h01;
		16'h8CED: out_word = 8'hC9;
		16'h8CEE: out_word = 8'hCD;
		16'h8CEF: out_word = 8'h1D;
		16'h8CF0: out_word = 8'h0B;
		16'h8CF1: out_word = 8'h79;
		16'h8CF2: out_word = 8'hCD;
		16'h8CF3: out_word = 8'hA3;
		16'h8CF4: out_word = 8'h11;
		16'h8CF5: out_word = 8'hC9;
		16'h8CF6: out_word = 8'hFD;
		16'h8CF7: out_word = 8'h36;
		16'h8CF8: out_word = 8'h10;
		16'h8CF9: out_word = 8'hFF;
		16'h8CFA: out_word = 8'hC9;
		16'h8CFB: out_word = 8'hCD;
		16'h8CFC: out_word = 8'h19;
		16'h8CFD: out_word = 8'h0E;
		16'h8CFE: out_word = 8'hDA;
		16'h8CFF: out_word = 8'h81;
		16'h8D00: out_word = 8'h0D;
		16'h8D01: out_word = 8'hCD;
		16'h8D02: out_word = 8'hAC;
		16'h8D03: out_word = 8'h0D;
		16'h8D04: out_word = 8'hCD;
		16'h8D05: out_word = 8'hB4;
		16'h8D06: out_word = 8'h0D;
		16'h8D07: out_word = 8'hAF;
		16'h8D08: out_word = 8'hDD;
		16'h8D09: out_word = 8'h77;
		16'h8D0A: out_word = 8'h21;
		16'h8D0B: out_word = 8'hCD;
		16'h8D0C: out_word = 8'hC8;
		16'h8D0D: out_word = 8'h0E;
		16'h8D0E: out_word = 8'hCD;
		16'h8D0F: out_word = 8'h1D;
		16'h8D10: out_word = 8'h0B;
		16'h8D11: out_word = 8'h79;
		16'h8D12: out_word = 8'hB7;
		16'h8D13: out_word = 8'hCA;
		16'h8D14: out_word = 8'h12;
		16'h8D15: out_word = 8'h0F;
		16'h8D16: out_word = 8'hFE;
		16'h8D17: out_word = 8'h0D;
		16'h8D18: out_word = 8'hD2;
		16'h8D19: out_word = 8'h12;
		16'h8D1A: out_word = 8'h0F;
		16'h8D1B: out_word = 8'hFE;
		16'h8D1C: out_word = 8'h0A;
		16'h8D1D: out_word = 8'h38;
		16'h8D1E: out_word = 8'h13;
		16'h8D1F: out_word = 8'hCD;
		16'h8D20: out_word = 8'h00;
		16'h8D21: out_word = 8'h0E;
		16'h8D22: out_word = 8'hCD;
		16'h8D23: out_word = 8'h74;
		16'h8D24: out_word = 8'h0D;
		16'h8D25: out_word = 8'h73;
		16'h8D26: out_word = 8'h23;
		16'h8D27: out_word = 8'h72;
		16'h8D28: out_word = 8'hCD;
		16'h8D29: out_word = 8'h74;
		16'h8D2A: out_word = 8'h0D;
		16'h8D2B: out_word = 8'h23;
		16'h8D2C: out_word = 8'h73;
		16'h8D2D: out_word = 8'h23;
		16'h8D2E: out_word = 8'h72;
		16'h8D2F: out_word = 8'h23;
		16'h8D30: out_word = 8'h18;
		16'h8D31: out_word = 8'h06;
		16'h8D32: out_word = 8'hDD;
		16'h8D33: out_word = 8'h71;
		16'h8D34: out_word = 8'h05;
		16'h8D35: out_word = 8'hCD;
		16'h8D36: out_word = 8'h00;
		16'h8D37: out_word = 8'h0E;
		16'h8D38: out_word = 8'hCD;
		16'h8D39: out_word = 8'h74;
		16'h8D3A: out_word = 8'h0D;
		16'h8D3B: out_word = 8'hCD;
		16'h8D3C: out_word = 8'hE3;
		16'h8D3D: out_word = 8'h0E;
		16'h8D3E: out_word = 8'hFE;
		16'h8D3F: out_word = 8'h5F;
		16'h8D40: out_word = 8'h20;
		16'h8D41: out_word = 8'h2C;
		16'h8D42: out_word = 8'hCD;
		16'h8D43: out_word = 8'hC5;
		16'h8D44: out_word = 8'h0A;
		16'h8D45: out_word = 8'hCD;
		16'h8D46: out_word = 8'h1D;
		16'h8D47: out_word = 8'h0B;
		16'h8D48: out_word = 8'h79;
		16'h8D49: out_word = 8'hFE;
		16'h8D4A: out_word = 8'h0A;
		16'h8D4B: out_word = 8'h38;
		16'h8D4C: out_word = 8'h12;
		16'h8D4D: out_word = 8'hE5;
		16'h8D4E: out_word = 8'hD5;
		16'h8D4F: out_word = 8'hCD;
		16'h8D50: out_word = 8'h00;
		16'h8D51: out_word = 8'h0E;
		16'h8D52: out_word = 8'hE1;
		16'h8D53: out_word = 8'h19;
		16'h8D54: out_word = 8'h4B;
		16'h8D55: out_word = 8'h42;
		16'h8D56: out_word = 8'hEB;
		16'h8D57: out_word = 8'hE1;
		16'h8D58: out_word = 8'h73;
		16'h8D59: out_word = 8'h23;
		16'h8D5A: out_word = 8'h72;
		16'h8D5B: out_word = 8'h59;
		16'h8D5C: out_word = 8'h50;
		16'h8D5D: out_word = 8'h18;
		16'h8D5E: out_word = 8'hC9;
		16'h8D5F: out_word = 8'hDD;
		16'h8D60: out_word = 8'h71;
		16'h8D61: out_word = 8'h05;
		16'h8D62: out_word = 8'hE5;
		16'h8D63: out_word = 8'hD5;
		16'h8D64: out_word = 8'hCD;
		16'h8D65: out_word = 8'h00;
		16'h8D66: out_word = 8'h0E;
		16'h8D67: out_word = 8'hE1;
		16'h8D68: out_word = 8'h19;
		16'h8D69: out_word = 8'hEB;
		16'h8D6A: out_word = 8'hE1;
		16'h8D6B: out_word = 8'hC3;
		16'h8D6C: out_word = 8'h3B;
		16'h8D6D: out_word = 8'h0D;
		16'h8D6E: out_word = 8'h73;
		16'h8D6F: out_word = 8'h23;
		16'h8D70: out_word = 8'h72;
		16'h8D71: out_word = 8'hC3;
		16'h8D72: out_word = 8'h9C;
		16'h8D73: out_word = 8'h0D;
		16'h8D74: out_word = 8'hDD;
		16'h8D75: out_word = 8'h7E;
		16'h8D76: out_word = 8'h21;
		16'h8D77: out_word = 8'h3C;
		16'h8D78: out_word = 8'hFE;
		16'h8D79: out_word = 8'h0B;
		16'h8D7A: out_word = 8'hCA;
		16'h8D7B: out_word = 8'h3A;
		16'h8D7C: out_word = 8'h0F;
		16'h8D7D: out_word = 8'hDD;
		16'h8D7E: out_word = 8'h77;
		16'h8D7F: out_word = 8'h21;
		16'h8D80: out_word = 8'hC9;
		16'h8D81: out_word = 8'hCD;
		16'h8D82: out_word = 8'hC8;
		16'h8D83: out_word = 8'h0E;
		16'h8D84: out_word = 8'hDD;
		16'h8D85: out_word = 8'h36;
		16'h8D86: out_word = 8'h21;
		16'h8D87: out_word = 8'h01;
		16'h8D88: out_word = 8'hCD;
		16'h8D89: out_word = 8'hAC;
		16'h8D8A: out_word = 8'h0D;
		16'h8D8B: out_word = 8'hCD;
		16'h8D8C: out_word = 8'hB4;
		16'h8D8D: out_word = 8'h0D;
		16'h8D8E: out_word = 8'hDD;
		16'h8D8F: out_word = 8'h4E;
		16'h8D90: out_word = 8'h05;
		16'h8D91: out_word = 8'hE5;
		16'h8D92: out_word = 8'hCD;
		16'h8D93: out_word = 8'h00;
		16'h8D94: out_word = 8'h0E;
		16'h8D95: out_word = 8'hE1;
		16'h8D96: out_word = 8'h73;
		16'h8D97: out_word = 8'h23;
		16'h8D98: out_word = 8'h72;
		16'h8D99: out_word = 8'hC3;
		16'h8D9A: out_word = 8'h9C;
		16'h8D9B: out_word = 8'h0D;
		16'h8D9C: out_word = 8'hE1;
		16'h8D9D: out_word = 8'h23;
		16'h8D9E: out_word = 8'h23;
		16'h8D9F: out_word = 8'hE5;
		16'h8DA0: out_word = 8'hC9;
		16'h8DA1: out_word = 8'hE1;
		16'h8DA2: out_word = 8'hFD;
		16'h8DA3: out_word = 8'h7E;
		16'h8DA4: out_word = 8'h21;
		16'h8DA5: out_word = 8'hFD;
		16'h8DA6: out_word = 8'hB6;
		16'h8DA7: out_word = 8'h10;
		16'h8DA8: out_word = 8'hFD;
		16'h8DA9: out_word = 8'h77;
		16'h8DAA: out_word = 8'h10;
		16'h8DAB: out_word = 8'hC9;
		16'h8DAC: out_word = 8'hDD;
		16'h8DAD: out_word = 8'hE5;
		16'h8DAE: out_word = 8'hE1;
		16'h8DAF: out_word = 8'h01;
		16'h8DB0: out_word = 8'h22;
		16'h8DB1: out_word = 8'h00;
		16'h8DB2: out_word = 8'h09;
		16'h8DB3: out_word = 8'hC9;
		16'h8DB4: out_word = 8'hE5;
		16'h8DB5: out_word = 8'hFD;
		16'h8DB6: out_word = 8'hE5;
		16'h8DB7: out_word = 8'hE1;
		16'h8DB8: out_word = 8'h01;
		16'h8DB9: out_word = 8'h11;
		16'h8DBA: out_word = 8'h00;
		16'h8DBB: out_word = 8'h09;
		16'h8DBC: out_word = 8'h06;
		16'h8DBD: out_word = 8'h00;
		16'h8DBE: out_word = 8'hDD;
		16'h8DBF: out_word = 8'h4E;
		16'h8DC0: out_word = 8'h02;
		16'h8DC1: out_word = 8'hCB;
		16'h8DC2: out_word = 8'h21;
		16'h8DC3: out_word = 8'h09;
		16'h8DC4: out_word = 8'hD1;
		16'h8DC5: out_word = 8'h73;
		16'h8DC6: out_word = 8'h23;
		16'h8DC7: out_word = 8'h72;
		16'h8DC8: out_word = 8'hEB;
		16'h8DC9: out_word = 8'hC9;
		16'h8DCA: out_word = 8'hFB;
		16'h8DCB: out_word = 8'h0C;
		16'h8DCC: out_word = 8'h85;
		16'h8DCD: out_word = 8'h0B;
		16'h8DCE: out_word = 8'h90;
		16'h8DCF: out_word = 8'h0B;
		16'h8DD0: out_word = 8'hA5;
		16'h8DD1: out_word = 8'h0B;
		16'h8DD2: out_word = 8'hA6;
		16'h8DD3: out_word = 8'h0B;
		16'h8DD4: out_word = 8'hC2;
		16'h8DD5: out_word = 8'h0B;
		16'h8DD6: out_word = 8'h32;
		16'h8DD7: out_word = 8'h0C;
		16'h8DD8: out_word = 8'h84;
		16'h8DD9: out_word = 8'h0C;
		16'h8DDA: out_word = 8'h95;
		16'h8DDB: out_word = 8'h0C;
		16'h8DDC: out_word = 8'hAD;
		16'h8DDD: out_word = 8'h0C;
		16'h8DDE: out_word = 8'hBA;
		16'h8DDF: out_word = 8'h0C;
		16'h8DE0: out_word = 8'hCE;
		16'h8DE1: out_word = 8'h0C;
		16'h8DE2: out_word = 8'hDD;
		16'h8DE3: out_word = 8'h0C;
		16'h8DE4: out_word = 8'hEE;
		16'h8DE5: out_word = 8'h0C;
		16'h8DE6: out_word = 8'hF6;
		16'h8DE7: out_word = 8'h0C;
		16'h8DE8: out_word = 8'h00;
		16'h8DE9: out_word = 8'h04;
		16'h8DEA: out_word = 8'h0B;
		16'h8DEB: out_word = 8'h0D;
		16'h8DEC: out_word = 8'h08;
		16'h8DED: out_word = 8'h0C;
		16'h8DEE: out_word = 8'h0E;
		16'h8DEF: out_word = 8'h0A;
		16'h8DF0: out_word = 8'h01;
		16'h8DF1: out_word = 8'h0F;
		16'h8DF2: out_word = 8'h00;
		16'h8DF3: out_word = 8'h21;
		16'h8DF4: out_word = 8'hB7;
		16'h8DF5: out_word = 8'h0A;
		16'h8DF6: out_word = 8'hED;
		16'h8DF7: out_word = 8'hB1;
		16'h8DF8: out_word = 8'hC9;
		16'h8DF9: out_word = 8'h09;
		16'h8DFA: out_word = 8'h0B;
		16'h8DFB: out_word = 8'h00;
		16'h8DFC: out_word = 8'h02;
		16'h8DFD: out_word = 8'h04;
		16'h8DFE: out_word = 8'h05;
		16'h8DFF: out_word = 8'h07;
		16'h8E00: out_word = 8'hE5;
		16'h8E01: out_word = 8'h06;
		16'h8E02: out_word = 8'h00;
		16'h8E03: out_word = 8'h21;
		16'h8E04: out_word = 8'h0C;
		16'h8E05: out_word = 8'h0E;
		16'h8E06: out_word = 8'h09;
		16'h8E07: out_word = 8'h16;
		16'h8E08: out_word = 8'h00;
		16'h8E09: out_word = 8'h5E;
		16'h8E0A: out_word = 8'hE1;
		16'h8E0B: out_word = 8'hC9;
		16'h8E0C: out_word = 8'h80;
		16'h8E0D: out_word = 8'h06;
		16'h8E0E: out_word = 8'h09;
		16'h8E0F: out_word = 8'h0C;
		16'h8E10: out_word = 8'h12;
		16'h8E11: out_word = 8'h18;
		16'h8E12: out_word = 8'h24;
		16'h8E13: out_word = 8'h30;
		16'h8E14: out_word = 8'h48;
		16'h8E15: out_word = 8'h60;
		16'h8E16: out_word = 8'h04;
		16'h8E17: out_word = 8'h08;
		16'h8E18: out_word = 8'h10;
		16'h8E19: out_word = 8'hFE;
		16'h8E1A: out_word = 8'h30;
		16'h8E1B: out_word = 8'hD8;
		16'h8E1C: out_word = 8'hFE;
		16'h8E1D: out_word = 8'h3A;
		16'h8E1E: out_word = 8'h3F;
		16'h8E1F: out_word = 8'hC9;
		16'h8E20: out_word = 8'h4F;
		16'h8E21: out_word = 8'hDD;
		16'h8E22: out_word = 8'h7E;
		16'h8E23: out_word = 8'h03;
		16'h8E24: out_word = 8'h81;
		16'h8E25: out_word = 8'hFE;
		16'h8E26: out_word = 8'h80;
		16'h8E27: out_word = 8'hD2;
		16'h8E28: out_word = 8'h32;
		16'h8E29: out_word = 8'h0F;
		16'h8E2A: out_word = 8'h4F;
		16'h8E2B: out_word = 8'hDD;
		16'h8E2C: out_word = 8'h7E;
		16'h8E2D: out_word = 8'h02;
		16'h8E2E: out_word = 8'hB7;
		16'h8E2F: out_word = 8'h20;
		16'h8E30: out_word = 8'h0E;
		16'h8E31: out_word = 8'h79;
		16'h8E32: out_word = 8'h2F;
		16'h8E33: out_word = 8'hE6;
		16'h8E34: out_word = 8'h7F;
		16'h8E35: out_word = 8'hCB;
		16'h8E36: out_word = 8'h3F;
		16'h8E37: out_word = 8'hCB;
		16'h8E38: out_word = 8'h3F;
		16'h8E39: out_word = 8'h16;
		16'h8E3A: out_word = 8'h06;
		16'h8E3B: out_word = 8'h5F;
		16'h8E3C: out_word = 8'hCD;
		16'h8E3D: out_word = 8'h7C;
		16'h8E3E: out_word = 8'h0E;
		16'h8E3F: out_word = 8'hDD;
		16'h8E40: out_word = 8'h71;
		16'h8E41: out_word = 8'h00;
		16'h8E42: out_word = 8'hDD;
		16'h8E43: out_word = 8'h7E;
		16'h8E44: out_word = 8'h02;
		16'h8E45: out_word = 8'hFE;
		16'h8E46: out_word = 8'h03;
		16'h8E47: out_word = 8'hD0;
		16'h8E48: out_word = 8'h21;
		16'h8E49: out_word = 8'h96;
		16'h8E4A: out_word = 8'h10;
		16'h8E4B: out_word = 8'h06;
		16'h8E4C: out_word = 8'h00;
		16'h8E4D: out_word = 8'h79;
		16'h8E4E: out_word = 8'hD6;
		16'h8E4F: out_word = 8'h15;
		16'h8E50: out_word = 8'h30;
		16'h8E51: out_word = 8'h05;
		16'h8E52: out_word = 8'h11;
		16'h8E53: out_word = 8'hBF;
		16'h8E54: out_word = 8'h0F;
		16'h8E55: out_word = 8'h18;
		16'h8E56: out_word = 8'h07;
		16'h8E57: out_word = 8'h4F;
		16'h8E58: out_word = 8'hCB;
		16'h8E59: out_word = 8'h21;
		16'h8E5A: out_word = 8'h09;
		16'h8E5B: out_word = 8'h5E;
		16'h8E5C: out_word = 8'h23;
		16'h8E5D: out_word = 8'h56;
		16'h8E5E: out_word = 8'hEB;
		16'h8E5F: out_word = 8'hDD;
		16'h8E60: out_word = 8'h56;
		16'h8E61: out_word = 8'h02;
		16'h8E62: out_word = 8'hCB;
		16'h8E63: out_word = 8'h22;
		16'h8E64: out_word = 8'h5D;
		16'h8E65: out_word = 8'hCD;
		16'h8E66: out_word = 8'h7C;
		16'h8E67: out_word = 8'h0E;
		16'h8E68: out_word = 8'h14;
		16'h8E69: out_word = 8'h5C;
		16'h8E6A: out_word = 8'hCD;
		16'h8E6B: out_word = 8'h7C;
		16'h8E6C: out_word = 8'h0E;
		16'h8E6D: out_word = 8'hDD;
		16'h8E6E: out_word = 8'hCB;
		16'h8E6F: out_word = 8'h04;
		16'h8E70: out_word = 8'h66;
		16'h8E71: out_word = 8'hC8;
		16'h8E72: out_word = 8'h16;
		16'h8E73: out_word = 8'h0D;
		16'h8E74: out_word = 8'hFD;
		16'h8E75: out_word = 8'h7E;
		16'h8E76: out_word = 8'h29;
		16'h8E77: out_word = 8'h5F;
		16'h8E78: out_word = 8'hCD;
		16'h8E79: out_word = 8'h7C;
		16'h8E7A: out_word = 8'h0E;
		16'h8E7B: out_word = 8'hC9;
		16'h8E7C: out_word = 8'hC5;
		16'h8E7D: out_word = 8'h01;
		16'h8E7E: out_word = 8'hFD;
		16'h8E7F: out_word = 8'hFF;
		16'h8E80: out_word = 8'hED;
		16'h8E81: out_word = 8'h51;
		16'h8E82: out_word = 8'h01;
		16'h8E83: out_word = 8'hFD;
		16'h8E84: out_word = 8'hBF;
		16'h8E85: out_word = 8'hED;
		16'h8E86: out_word = 8'h59;
		16'h8E87: out_word = 8'hC1;
		16'h8E88: out_word = 8'hC9;
		16'h8E89: out_word = 8'hC5;
		16'h8E8A: out_word = 8'h01;
		16'h8E8B: out_word = 8'hFD;
		16'h8E8C: out_word = 8'hFF;
		16'h8E8D: out_word = 8'hED;
		16'h8E8E: out_word = 8'h79;
		16'h8E8F: out_word = 8'hED;
		16'h8E90: out_word = 8'h78;
		16'h8E91: out_word = 8'hC1;
		16'h8E92: out_word = 8'hC9;
		16'h8E93: out_word = 8'h16;
		16'h8E94: out_word = 8'h07;
		16'h8E95: out_word = 8'h1E;
		16'h8E96: out_word = 8'hFF;
		16'h8E97: out_word = 8'hCD;
		16'h8E98: out_word = 8'h7C;
		16'h8E99: out_word = 8'h0E;
		16'h8E9A: out_word = 8'h16;
		16'h8E9B: out_word = 8'h08;
		16'h8E9C: out_word = 8'h1E;
		16'h8E9D: out_word = 8'h00;
		16'h8E9E: out_word = 8'hCD;
		16'h8E9F: out_word = 8'h7C;
		16'h8EA0: out_word = 8'h0E;
		16'h8EA1: out_word = 8'h14;
		16'h8EA2: out_word = 8'hCD;
		16'h8EA3: out_word = 8'h7C;
		16'h8EA4: out_word = 8'h0E;
		16'h8EA5: out_word = 8'h14;
		16'h8EA6: out_word = 8'hCD;
		16'h8EA7: out_word = 8'h7C;
		16'h8EA8: out_word = 8'h0E;
		16'h8EA9: out_word = 8'hCD;
		16'h8EAA: out_word = 8'h4F;
		16'h8EAB: out_word = 8'h0A;
		16'h8EAC: out_word = 8'hFD;
		16'h8EAD: out_word = 8'hCB;
		16'h8EAE: out_word = 8'h22;
		16'h8EAF: out_word = 8'h1E;
		16'h8EB0: out_word = 8'h38;
		16'h8EB1: out_word = 8'h06;
		16'h8EB2: out_word = 8'hCD;
		16'h8EB3: out_word = 8'h67;
		16'h8EB4: out_word = 8'h0A;
		16'h8EB5: out_word = 8'hCD;
		16'h8EB6: out_word = 8'h8D;
		16'h8EB7: out_word = 8'h11;
		16'h8EB8: out_word = 8'hFD;
		16'h8EB9: out_word = 8'hCB;
		16'h8EBA: out_word = 8'h21;
		16'h8EBB: out_word = 8'h26;
		16'h8EBC: out_word = 8'h38;
		16'h8EBD: out_word = 8'h05;
		16'h8EBE: out_word = 8'hCD;
		16'h8EBF: out_word = 8'h6E;
		16'h8EC0: out_word = 8'h0A;
		16'h8EC1: out_word = 8'h18;
		16'h8EC2: out_word = 8'hE9;
		16'h8EC3: out_word = 8'hFD;
		16'h8EC4: out_word = 8'h21;
		16'h8EC5: out_word = 8'h3A;
		16'h8EC6: out_word = 8'h5C;
		16'h8EC7: out_word = 8'hC9;
		16'h8EC8: out_word = 8'hE5;
		16'h8EC9: out_word = 8'hD5;
		16'h8ECA: out_word = 8'hDD;
		16'h8ECB: out_word = 8'h6E;
		16'h8ECC: out_word = 8'h06;
		16'h8ECD: out_word = 8'hDD;
		16'h8ECE: out_word = 8'h66;
		16'h8ECF: out_word = 8'h07;
		16'h8ED0: out_word = 8'h2B;
		16'h8ED1: out_word = 8'h7E;
		16'h8ED2: out_word = 8'hFE;
		16'h8ED3: out_word = 8'h20;
		16'h8ED4: out_word = 8'h28;
		16'h8ED5: out_word = 8'hFA;
		16'h8ED6: out_word = 8'hFE;
		16'h8ED7: out_word = 8'h0D;
		16'h8ED8: out_word = 8'h28;
		16'h8ED9: out_word = 8'hF6;
		16'h8EDA: out_word = 8'hDD;
		16'h8EDB: out_word = 8'h75;
		16'h8EDC: out_word = 8'h06;
		16'h8EDD: out_word = 8'hDD;
		16'h8EDE: out_word = 8'h74;
		16'h8EDF: out_word = 8'h07;
		16'h8EE0: out_word = 8'hD1;
		16'h8EE1: out_word = 8'hE1;
		16'h8EE2: out_word = 8'hC9;
		16'h8EE3: out_word = 8'hE5;
		16'h8EE4: out_word = 8'hD5;
		16'h8EE5: out_word = 8'hC5;
		16'h8EE6: out_word = 8'hDD;
		16'h8EE7: out_word = 8'h6E;
		16'h8EE8: out_word = 8'h06;
		16'h8EE9: out_word = 8'hDD;
		16'h8EEA: out_word = 8'h66;
		16'h8EEB: out_word = 8'h07;
		16'h8EEC: out_word = 8'h7C;
		16'h8EED: out_word = 8'hDD;
		16'h8EEE: out_word = 8'hBE;
		16'h8EEF: out_word = 8'h09;
		16'h8EF0: out_word = 8'h20;
		16'h8EF1: out_word = 8'h09;
		16'h8EF2: out_word = 8'h7D;
		16'h8EF3: out_word = 8'hDD;
		16'h8EF4: out_word = 8'hBE;
		16'h8EF5: out_word = 8'h08;
		16'h8EF6: out_word = 8'h20;
		16'h8EF7: out_word = 8'h03;
		16'h8EF8: out_word = 8'h37;
		16'h8EF9: out_word = 8'h18;
		16'h8EFA: out_word = 8'h0A;
		16'h8EFB: out_word = 8'h7E;
		16'h8EFC: out_word = 8'hFE;
		16'h8EFD: out_word = 8'h20;
		16'h8EFE: out_word = 8'h28;
		16'h8EFF: out_word = 8'h09;
		16'h8F00: out_word = 8'hFE;
		16'h8F01: out_word = 8'h0D;
		16'h8F02: out_word = 8'h28;
		16'h8F03: out_word = 8'h05;
		16'h8F04: out_word = 8'hB7;
		16'h8F05: out_word = 8'hC1;
		16'h8F06: out_word = 8'hD1;
		16'h8F07: out_word = 8'hE1;
		16'h8F08: out_word = 8'hC9;
		16'h8F09: out_word = 8'h23;
		16'h8F0A: out_word = 8'hDD;
		16'h8F0B: out_word = 8'h75;
		16'h8F0C: out_word = 8'h06;
		16'h8F0D: out_word = 8'hDD;
		16'h8F0E: out_word = 8'h74;
		16'h8F0F: out_word = 8'h07;
		16'h8F10: out_word = 8'h18;
		16'h8F11: out_word = 8'hDA;
		16'h8F12: out_word = 8'hCD;
		16'h8F13: out_word = 8'h93;
		16'h8F14: out_word = 8'h0E;
		16'h8F15: out_word = 8'hFB;
		16'h8F16: out_word = 8'hCD;
		16'h8F17: out_word = 8'hAC;
		16'h8F18: out_word = 8'h05;
		16'h8F19: out_word = 8'h29;
		16'h8F1A: out_word = 8'hCD;
		16'h8F1B: out_word = 8'h93;
		16'h8F1C: out_word = 8'h0E;
		16'h8F1D: out_word = 8'hFB;
		16'h8F1E: out_word = 8'hCD;
		16'h8F1F: out_word = 8'hAC;
		16'h8F20: out_word = 8'h05;
		16'h8F21: out_word = 8'h27;
		16'h8F22: out_word = 8'hCD;
		16'h8F23: out_word = 8'h93;
		16'h8F24: out_word = 8'h0E;
		16'h8F25: out_word = 8'hFB;
		16'h8F26: out_word = 8'hCD;
		16'h8F27: out_word = 8'hAC;
		16'h8F28: out_word = 8'h05;
		16'h8F29: out_word = 8'h26;
		16'h8F2A: out_word = 8'hCD;
		16'h8F2B: out_word = 8'h93;
		16'h8F2C: out_word = 8'h0E;
		16'h8F2D: out_word = 8'hFB;
		16'h8F2E: out_word = 8'hCD;
		16'h8F2F: out_word = 8'hAC;
		16'h8F30: out_word = 8'h05;
		16'h8F31: out_word = 8'h1F;
		16'h8F32: out_word = 8'hCD;
		16'h8F33: out_word = 8'h93;
		16'h8F34: out_word = 8'h0E;
		16'h8F35: out_word = 8'hFB;
		16'h8F36: out_word = 8'hCD;
		16'h8F37: out_word = 8'hAC;
		16'h8F38: out_word = 8'h05;
		16'h8F39: out_word = 8'h28;
		16'h8F3A: out_word = 8'hCD;
		16'h8F3B: out_word = 8'h93;
		16'h8F3C: out_word = 8'h0E;
		16'h8F3D: out_word = 8'hFB;
		16'h8F3E: out_word = 8'hCD;
		16'h8F3F: out_word = 8'hAC;
		16'h8F40: out_word = 8'h05;
		16'h8F41: out_word = 8'h2A;
		16'h8F42: out_word = 8'hCD;
		16'h8F43: out_word = 8'h4F;
		16'h8F44: out_word = 8'h0A;
		16'h8F45: out_word = 8'hFD;
		16'h8F46: out_word = 8'hCB;
		16'h8F47: out_word = 8'h22;
		16'h8F48: out_word = 8'h1E;
		16'h8F49: out_word = 8'h38;
		16'h8F4A: out_word = 8'h21;
		16'h8F4B: out_word = 8'hCD;
		16'h8F4C: out_word = 8'h67;
		16'h8F4D: out_word = 8'h0A;
		16'h8F4E: out_word = 8'hCD;
		16'h8F4F: out_word = 8'hD1;
		16'h8F50: out_word = 8'h0A;
		16'h8F51: out_word = 8'hFE;
		16'h8F52: out_word = 8'h80;
		16'h8F53: out_word = 8'h28;
		16'h8F54: out_word = 8'h17;
		16'h8F55: out_word = 8'hCD;
		16'h8F56: out_word = 8'h20;
		16'h8F57: out_word = 8'h0E;
		16'h8F58: out_word = 8'hDD;
		16'h8F59: out_word = 8'h7E;
		16'h8F5A: out_word = 8'h02;
		16'h8F5B: out_word = 8'hFE;
		16'h8F5C: out_word = 8'h03;
		16'h8F5D: out_word = 8'h30;
		16'h8F5E: out_word = 8'h0A;
		16'h8F5F: out_word = 8'h16;
		16'h8F60: out_word = 8'h08;
		16'h8F61: out_word = 8'h82;
		16'h8F62: out_word = 8'h57;
		16'h8F63: out_word = 8'hDD;
		16'h8F64: out_word = 8'h5E;
		16'h8F65: out_word = 8'h04;
		16'h8F66: out_word = 8'hCD;
		16'h8F67: out_word = 8'h7C;
		16'h8F68: out_word = 8'h0E;
		16'h8F69: out_word = 8'hCD;
		16'h8F6A: out_word = 8'h6E;
		16'h8F6B: out_word = 8'h11;
		16'h8F6C: out_word = 8'hFD;
		16'h8F6D: out_word = 8'hCB;
		16'h8F6E: out_word = 8'h21;
		16'h8F6F: out_word = 8'h26;
		16'h8F70: out_word = 8'hD8;
		16'h8F71: out_word = 8'hCD;
		16'h8F72: out_word = 8'h6E;
		16'h8F73: out_word = 8'h0A;
		16'h8F74: out_word = 8'h18;
		16'h8F75: out_word = 8'hCF;
		16'h8F76: out_word = 8'hE5;
		16'h8F77: out_word = 8'hFD;
		16'h8F78: out_word = 8'h6E;
		16'h8F79: out_word = 8'h27;
		16'h8F7A: out_word = 8'hFD;
		16'h8F7B: out_word = 8'h66;
		16'h8F7C: out_word = 8'h28;
		16'h8F7D: out_word = 8'h01;
		16'h8F7E: out_word = 8'h64;
		16'h8F7F: out_word = 8'h00;
		16'h8F80: out_word = 8'hB7;
		16'h8F81: out_word = 8'hED;
		16'h8F82: out_word = 8'h42;
		16'h8F83: out_word = 8'hE5;
		16'h8F84: out_word = 8'hC1;
		16'h8F85: out_word = 8'hE1;
		16'h8F86: out_word = 8'h0B;
		16'h8F87: out_word = 8'h78;
		16'h8F88: out_word = 8'hB1;
		16'h8F89: out_word = 8'h20;
		16'h8F8A: out_word = 8'hFB;
		16'h8F8B: out_word = 8'h1B;
		16'h8F8C: out_word = 8'h7A;
		16'h8F8D: out_word = 8'hB3;
		16'h8F8E: out_word = 8'h20;
		16'h8F8F: out_word = 8'hE6;
		16'h8F90: out_word = 8'hC9;
		16'h8F91: out_word = 8'h11;
		16'h8F92: out_word = 8'hFF;
		16'h8F93: out_word = 8'hFF;
		16'h8F94: out_word = 8'hCD;
		16'h8F95: out_word = 8'h4A;
		16'h8F96: out_word = 8'h0A;
		16'h8F97: out_word = 8'hFD;
		16'h8F98: out_word = 8'hCB;
		16'h8F99: out_word = 8'h22;
		16'h8F9A: out_word = 8'h1E;
		16'h8F9B: out_word = 8'h38;
		16'h8F9C: out_word = 8'h12;
		16'h8F9D: out_word = 8'hD5;
		16'h8F9E: out_word = 8'h5E;
		16'h8F9F: out_word = 8'h23;
		16'h8FA0: out_word = 8'h56;
		16'h8FA1: out_word = 8'hEB;
		16'h8FA2: out_word = 8'h5E;
		16'h8FA3: out_word = 8'h23;
		16'h8FA4: out_word = 8'h56;
		16'h8FA5: out_word = 8'hD5;
		16'h8FA6: out_word = 8'hE1;
		16'h8FA7: out_word = 8'hC1;
		16'h8FA8: out_word = 8'hB7;
		16'h8FA9: out_word = 8'hED;
		16'h8FAA: out_word = 8'h42;
		16'h8FAB: out_word = 8'h38;
		16'h8FAC: out_word = 8'h02;
		16'h8FAD: out_word = 8'hC5;
		16'h8FAE: out_word = 8'hD1;
		16'h8FAF: out_word = 8'hFD;
		16'h8FB0: out_word = 8'hCB;
		16'h8FB1: out_word = 8'h21;
		16'h8FB2: out_word = 8'h26;
		16'h8FB3: out_word = 8'h38;
		16'h8FB4: out_word = 8'h05;
		16'h8FB5: out_word = 8'hCD;
		16'h8FB6: out_word = 8'h6E;
		16'h8FB7: out_word = 8'h0A;
		16'h8FB8: out_word = 8'h18;
		16'h8FB9: out_word = 8'hDD;
		16'h8FBA: out_word = 8'hFD;
		16'h8FBB: out_word = 8'h73;
		16'h8FBC: out_word = 8'h25;
		16'h8FBD: out_word = 8'hFD;
		16'h8FBE: out_word = 8'h72;
		16'h8FBF: out_word = 8'h26;
		16'h8FC0: out_word = 8'hC9;
		16'h8FC1: out_word = 8'hAF;
		16'h8FC2: out_word = 8'hFD;
		16'h8FC3: out_word = 8'h77;
		16'h8FC4: out_word = 8'h2A;
		16'h8FC5: out_word = 8'hCD;
		16'h8FC6: out_word = 8'h4F;
		16'h8FC7: out_word = 8'h0A;
		16'h8FC8: out_word = 8'hFD;
		16'h8FC9: out_word = 8'hCB;
		16'h8FCA: out_word = 8'h22;
		16'h8FCB: out_word = 8'h1E;
		16'h8FCC: out_word = 8'hDA;
		16'h8FCD: out_word = 8'h5A;
		16'h8FCE: out_word = 8'h10;
		16'h8FCF: out_word = 8'hCD;
		16'h8FD0: out_word = 8'h67;
		16'h8FD1: out_word = 8'h0A;
		16'h8FD2: out_word = 8'hFD;
		16'h8FD3: out_word = 8'hE5;
		16'h8FD4: out_word = 8'hE1;
		16'h8FD5: out_word = 8'h01;
		16'h8FD6: out_word = 8'h11;
		16'h8FD7: out_word = 8'h00;
		16'h8FD8: out_word = 8'h09;
		16'h8FD9: out_word = 8'h06;
		16'h8FDA: out_word = 8'h00;
		16'h8FDB: out_word = 8'hDD;
		16'h8FDC: out_word = 8'h4E;
		16'h8FDD: out_word = 8'h02;
		16'h8FDE: out_word = 8'hCB;
		16'h8FDF: out_word = 8'h21;
		16'h8FE0: out_word = 8'h09;
		16'h8FE1: out_word = 8'h5E;
		16'h8FE2: out_word = 8'h23;
		16'h8FE3: out_word = 8'h56;
		16'h8FE4: out_word = 8'hEB;
		16'h8FE5: out_word = 8'hE5;
		16'h8FE6: out_word = 8'h5E;
		16'h8FE7: out_word = 8'h23;
		16'h8FE8: out_word = 8'h56;
		16'h8FE9: out_word = 8'hEB;
		16'h8FEA: out_word = 8'hFD;
		16'h8FEB: out_word = 8'h5E;
		16'h8FEC: out_word = 8'h25;
		16'h8FED: out_word = 8'hFD;
		16'h8FEE: out_word = 8'h56;
		16'h8FEF: out_word = 8'h26;
		16'h8FF0: out_word = 8'hB7;
		16'h8FF1: out_word = 8'hED;
		16'h8FF2: out_word = 8'h52;
		16'h8FF3: out_word = 8'hEB;
		16'h8FF4: out_word = 8'hE1;
		16'h8FF5: out_word = 8'h28;
		16'h8FF6: out_word = 8'h05;
		16'h8FF7: out_word = 8'h73;
		16'h8FF8: out_word = 8'h23;
		16'h8FF9: out_word = 8'h72;
		16'h8FFA: out_word = 8'h18;
		16'h8FFB: out_word = 8'h5E;
		16'h8FFC: out_word = 8'hDD;
		16'h8FFD: out_word = 8'h7E;
		16'h8FFE: out_word = 8'h02;
		16'h8FFF: out_word = 8'hFE;
		16'h9000: out_word = 8'h03;
		16'h9001: out_word = 8'h30;
		16'h9002: out_word = 8'h09;
		16'h9003: out_word = 8'h16;
		16'h9004: out_word = 8'h08;
		16'h9005: out_word = 8'h82;
		16'h9006: out_word = 8'h57;
		16'h9007: out_word = 8'h1E;
		16'h9008: out_word = 8'h00;
		16'h9009: out_word = 8'hCD;
		16'h900A: out_word = 8'h7C;
		16'h900B: out_word = 8'h0E;
		16'h900C: out_word = 8'hCD;
		16'h900D: out_word = 8'h8D;
		16'h900E: out_word = 8'h11;
		16'h900F: out_word = 8'hDD;
		16'h9010: out_word = 8'hE5;
		16'h9011: out_word = 8'hE1;
		16'h9012: out_word = 8'h01;
		16'h9013: out_word = 8'h21;
		16'h9014: out_word = 8'h00;
		16'h9015: out_word = 8'h09;
		16'h9016: out_word = 8'h35;
		16'h9017: out_word = 8'h20;
		16'h9018: out_word = 8'h0D;
		16'h9019: out_word = 8'hCD;
		16'h901A: out_word = 8'h5C;
		16'h901B: out_word = 8'h0B;
		16'h901C: out_word = 8'hFD;
		16'h901D: out_word = 8'h7E;
		16'h901E: out_word = 8'h21;
		16'h901F: out_word = 8'hFD;
		16'h9020: out_word = 8'hA6;
		16'h9021: out_word = 8'h10;
		16'h9022: out_word = 8'h20;
		16'h9023: out_word = 8'h36;
		16'h9024: out_word = 8'h18;
		16'h9025: out_word = 8'h17;
		16'h9026: out_word = 8'hFD;
		16'h9027: out_word = 8'hE5;
		16'h9028: out_word = 8'hE1;
		16'h9029: out_word = 8'h01;
		16'h902A: out_word = 8'h11;
		16'h902B: out_word = 8'h00;
		16'h902C: out_word = 8'h09;
		16'h902D: out_word = 8'h06;
		16'h902E: out_word = 8'h00;
		16'h902F: out_word = 8'hDD;
		16'h9030: out_word = 8'h4E;
		16'h9031: out_word = 8'h02;
		16'h9032: out_word = 8'hCB;
		16'h9033: out_word = 8'h21;
		16'h9034: out_word = 8'h09;
		16'h9035: out_word = 8'h5E;
		16'h9036: out_word = 8'h23;
		16'h9037: out_word = 8'h56;
		16'h9038: out_word = 8'h13;
		16'h9039: out_word = 8'h13;
		16'h903A: out_word = 8'h72;
		16'h903B: out_word = 8'h2B;
		16'h903C: out_word = 8'h73;
		16'h903D: out_word = 8'hCD;
		16'h903E: out_word = 8'hD1;
		16'h903F: out_word = 8'h0A;
		16'h9040: out_word = 8'h4F;
		16'h9041: out_word = 8'hFD;
		16'h9042: out_word = 8'h7E;
		16'h9043: out_word = 8'h21;
		16'h9044: out_word = 8'hFD;
		16'h9045: out_word = 8'hA6;
		16'h9046: out_word = 8'h10;
		16'h9047: out_word = 8'h20;
		16'h9048: out_word = 8'h11;
		16'h9049: out_word = 8'h79;
		16'h904A: out_word = 8'hFE;
		16'h904B: out_word = 8'h80;
		16'h904C: out_word = 8'h28;
		16'h904D: out_word = 8'h0C;
		16'h904E: out_word = 8'hCD;
		16'h904F: out_word = 8'h20;
		16'h9050: out_word = 8'h0E;
		16'h9051: out_word = 8'hFD;
		16'h9052: out_word = 8'h7E;
		16'h9053: out_word = 8'h21;
		16'h9054: out_word = 8'hFD;
		16'h9055: out_word = 8'hB6;
		16'h9056: out_word = 8'h2A;
		16'h9057: out_word = 8'hFD;
		16'h9058: out_word = 8'h77;
		16'h9059: out_word = 8'h2A;
		16'h905A: out_word = 8'hFD;
		16'h905B: out_word = 8'hCB;
		16'h905C: out_word = 8'h21;
		16'h905D: out_word = 8'h26;
		16'h905E: out_word = 8'h38;
		16'h905F: out_word = 8'h06;
		16'h9060: out_word = 8'hCD;
		16'h9061: out_word = 8'h6E;
		16'h9062: out_word = 8'h0A;
		16'h9063: out_word = 8'hC3;
		16'h9064: out_word = 8'hC8;
		16'h9065: out_word = 8'h0F;
		16'h9066: out_word = 8'h11;
		16'h9067: out_word = 8'h01;
		16'h9068: out_word = 8'h00;
		16'h9069: out_word = 8'hCD;
		16'h906A: out_word = 8'h76;
		16'h906B: out_word = 8'h0F;
		16'h906C: out_word = 8'hCD;
		16'h906D: out_word = 8'h4F;
		16'h906E: out_word = 8'h0A;
		16'h906F: out_word = 8'hFD;
		16'h9070: out_word = 8'hCB;
		16'h9071: out_word = 8'h2A;
		16'h9072: out_word = 8'h1E;
		16'h9073: out_word = 8'h30;
		16'h9074: out_word = 8'h17;
		16'h9075: out_word = 8'hCD;
		16'h9076: out_word = 8'h67;
		16'h9077: out_word = 8'h0A;
		16'h9078: out_word = 8'hDD;
		16'h9079: out_word = 8'h7E;
		16'h907A: out_word = 8'h02;
		16'h907B: out_word = 8'hFE;
		16'h907C: out_word = 8'h03;
		16'h907D: out_word = 8'h30;
		16'h907E: out_word = 8'h0A;
		16'h907F: out_word = 8'h16;
		16'h9080: out_word = 8'h08;
		16'h9081: out_word = 8'h82;
		16'h9082: out_word = 8'h57;
		16'h9083: out_word = 8'hDD;
		16'h9084: out_word = 8'h5E;
		16'h9085: out_word = 8'h04;
		16'h9086: out_word = 8'hCD;
		16'h9087: out_word = 8'h7C;
		16'h9088: out_word = 8'h0E;
		16'h9089: out_word = 8'hCD;
		16'h908A: out_word = 8'h6E;
		16'h908B: out_word = 8'h11;
		16'h908C: out_word = 8'hFD;
		16'h908D: out_word = 8'hCB;
		16'h908E: out_word = 8'h21;
		16'h908F: out_word = 8'h26;
		16'h9090: out_word = 8'hD8;
		16'h9091: out_word = 8'hCD;
		16'h9092: out_word = 8'h6E;
		16'h9093: out_word = 8'h0A;
		16'h9094: out_word = 8'h18;
		16'h9095: out_word = 8'hD9;
		16'h9096: out_word = 8'hBF;
		16'h9097: out_word = 8'h0F;
		16'h9098: out_word = 8'hDC;
		16'h9099: out_word = 8'h0E;
		16'h909A: out_word = 8'h07;
		16'h909B: out_word = 8'h0E;
		16'h909C: out_word = 8'h3D;
		16'h909D: out_word = 8'h0D;
		16'h909E: out_word = 8'h7F;
		16'h909F: out_word = 8'h0C;
		16'h90A0: out_word = 8'hCC;
		16'h90A1: out_word = 8'h0B;
		16'h90A2: out_word = 8'h22;
		16'h90A3: out_word = 8'h0B;
		16'h90A4: out_word = 8'h82;
		16'h90A5: out_word = 8'h0A;
		16'h90A6: out_word = 8'hEB;
		16'h90A7: out_word = 8'h09;
		16'h90A8: out_word = 8'h5D;
		16'h90A9: out_word = 8'h09;
		16'h90AA: out_word = 8'hD6;
		16'h90AB: out_word = 8'h08;
		16'h90AC: out_word = 8'h57;
		16'h90AD: out_word = 8'h08;
		16'h90AE: out_word = 8'hDF;
		16'h90AF: out_word = 8'h07;
		16'h90B0: out_word = 8'h6E;
		16'h90B1: out_word = 8'h07;
		16'h90B2: out_word = 8'h03;
		16'h90B3: out_word = 8'h07;
		16'h90B4: out_word = 8'h9F;
		16'h90B5: out_word = 8'h06;
		16'h90B6: out_word = 8'h40;
		16'h90B7: out_word = 8'h06;
		16'h90B8: out_word = 8'hE6;
		16'h90B9: out_word = 8'h05;
		16'h90BA: out_word = 8'h91;
		16'h90BB: out_word = 8'h05;
		16'h90BC: out_word = 8'h41;
		16'h90BD: out_word = 8'h05;
		16'h90BE: out_word = 8'hF6;
		16'h90BF: out_word = 8'h04;
		16'h90C0: out_word = 8'hAE;
		16'h90C1: out_word = 8'h04;
		16'h90C2: out_word = 8'h6B;
		16'h90C3: out_word = 8'h04;
		16'h90C4: out_word = 8'h2C;
		16'h90C5: out_word = 8'h04;
		16'h90C6: out_word = 8'hF0;
		16'h90C7: out_word = 8'h03;
		16'h90C8: out_word = 8'hB7;
		16'h90C9: out_word = 8'h03;
		16'h90CA: out_word = 8'h82;
		16'h90CB: out_word = 8'h03;
		16'h90CC: out_word = 8'h4F;
		16'h90CD: out_word = 8'h03;
		16'h90CE: out_word = 8'h20;
		16'h90CF: out_word = 8'h03;
		16'h90D0: out_word = 8'hF3;
		16'h90D1: out_word = 8'h02;
		16'h90D2: out_word = 8'hC8;
		16'h90D3: out_word = 8'h02;
		16'h90D4: out_word = 8'hA1;
		16'h90D5: out_word = 8'h02;
		16'h90D6: out_word = 8'h7B;
		16'h90D7: out_word = 8'h02;
		16'h90D8: out_word = 8'h57;
		16'h90D9: out_word = 8'h02;
		16'h90DA: out_word = 8'h36;
		16'h90DB: out_word = 8'h02;
		16'h90DC: out_word = 8'h16;
		16'h90DD: out_word = 8'h02;
		16'h90DE: out_word = 8'hF8;
		16'h90DF: out_word = 8'h01;
		16'h90E0: out_word = 8'hDC;
		16'h90E1: out_word = 8'h01;
		16'h90E2: out_word = 8'hC1;
		16'h90E3: out_word = 8'h01;
		16'h90E4: out_word = 8'hA8;
		16'h90E5: out_word = 8'h01;
		16'h90E6: out_word = 8'h90;
		16'h90E7: out_word = 8'h01;
		16'h90E8: out_word = 8'h79;
		16'h90E9: out_word = 8'h01;
		16'h90EA: out_word = 8'h64;
		16'h90EB: out_word = 8'h01;
		16'h90EC: out_word = 8'h50;
		16'h90ED: out_word = 8'h01;
		16'h90EE: out_word = 8'h3D;
		16'h90EF: out_word = 8'h01;
		16'h90F0: out_word = 8'h2C;
		16'h90F1: out_word = 8'h01;
		16'h90F2: out_word = 8'h1B;
		16'h90F3: out_word = 8'h01;
		16'h90F4: out_word = 8'h0B;
		16'h90F5: out_word = 8'h01;
		16'h90F6: out_word = 8'hFC;
		16'h90F7: out_word = 8'h00;
		16'h90F8: out_word = 8'hEE;
		16'h90F9: out_word = 8'h00;
		16'h90FA: out_word = 8'hE0;
		16'h90FB: out_word = 8'h00;
		16'h90FC: out_word = 8'hD4;
		16'h90FD: out_word = 8'h00;
		16'h90FE: out_word = 8'hC8;
		16'h90FF: out_word = 8'h00;
		16'h9100: out_word = 8'hBD;
		16'h9101: out_word = 8'h00;
		16'h9102: out_word = 8'hB2;
		16'h9103: out_word = 8'h00;
		16'h9104: out_word = 8'hA8;
		16'h9105: out_word = 8'h00;
		16'h9106: out_word = 8'h9F;
		16'h9107: out_word = 8'h00;
		16'h9108: out_word = 8'h96;
		16'h9109: out_word = 8'h00;
		16'h910A: out_word = 8'h8D;
		16'h910B: out_word = 8'h00;
		16'h910C: out_word = 8'h85;
		16'h910D: out_word = 8'h00;
		16'h910E: out_word = 8'h7E;
		16'h910F: out_word = 8'h00;
		16'h9110: out_word = 8'h77;
		16'h9111: out_word = 8'h00;
		16'h9112: out_word = 8'h70;
		16'h9113: out_word = 8'h00;
		16'h9114: out_word = 8'h6A;
		16'h9115: out_word = 8'h00;
		16'h9116: out_word = 8'h64;
		16'h9117: out_word = 8'h00;
		16'h9118: out_word = 8'h5E;
		16'h9119: out_word = 8'h00;
		16'h911A: out_word = 8'h59;
		16'h911B: out_word = 8'h00;
		16'h911C: out_word = 8'h54;
		16'h911D: out_word = 8'h00;
		16'h911E: out_word = 8'h4F;
		16'h911F: out_word = 8'h00;
		16'h9120: out_word = 8'h4B;
		16'h9121: out_word = 8'h00;
		16'h9122: out_word = 8'h47;
		16'h9123: out_word = 8'h00;
		16'h9124: out_word = 8'h43;
		16'h9125: out_word = 8'h00;
		16'h9126: out_word = 8'h3F;
		16'h9127: out_word = 8'h00;
		16'h9128: out_word = 8'h3B;
		16'h9129: out_word = 8'h00;
		16'h912A: out_word = 8'h38;
		16'h912B: out_word = 8'h00;
		16'h912C: out_word = 8'h35;
		16'h912D: out_word = 8'h00;
		16'h912E: out_word = 8'h32;
		16'h912F: out_word = 8'h00;
		16'h9130: out_word = 8'h2F;
		16'h9131: out_word = 8'h00;
		16'h9132: out_word = 8'h2D;
		16'h9133: out_word = 8'h00;
		16'h9134: out_word = 8'h2A;
		16'h9135: out_word = 8'h00;
		16'h9136: out_word = 8'h28;
		16'h9137: out_word = 8'h00;
		16'h9138: out_word = 8'h25;
		16'h9139: out_word = 8'h00;
		16'h913A: out_word = 8'h23;
		16'h913B: out_word = 8'h00;
		16'h913C: out_word = 8'h21;
		16'h913D: out_word = 8'h00;
		16'h913E: out_word = 8'h1F;
		16'h913F: out_word = 8'h00;
		16'h9140: out_word = 8'h1E;
		16'h9141: out_word = 8'h00;
		16'h9142: out_word = 8'h1C;
		16'h9143: out_word = 8'h00;
		16'h9144: out_word = 8'h1A;
		16'h9145: out_word = 8'h00;
		16'h9146: out_word = 8'h19;
		16'h9147: out_word = 8'h00;
		16'h9148: out_word = 8'h18;
		16'h9149: out_word = 8'h00;
		16'h914A: out_word = 8'h16;
		16'h914B: out_word = 8'h00;
		16'h914C: out_word = 8'h15;
		16'h914D: out_word = 8'h00;
		16'h914E: out_word = 8'h14;
		16'h914F: out_word = 8'h00;
		16'h9150: out_word = 8'h13;
		16'h9151: out_word = 8'h00;
		16'h9152: out_word = 8'h12;
		16'h9153: out_word = 8'h00;
		16'h9154: out_word = 8'h11;
		16'h9155: out_word = 8'h00;
		16'h9156: out_word = 8'h10;
		16'h9157: out_word = 8'h00;
		16'h9158: out_word = 8'h0F;
		16'h9159: out_word = 8'h00;
		16'h915A: out_word = 8'h0E;
		16'h915B: out_word = 8'h00;
		16'h915C: out_word = 8'h0D;
		16'h915D: out_word = 8'h00;
		16'h915E: out_word = 8'h0C;
		16'h915F: out_word = 8'h00;
		16'h9160: out_word = 8'h0C;
		16'h9161: out_word = 8'h00;
		16'h9162: out_word = 8'h0B;
		16'h9163: out_word = 8'h00;
		16'h9164: out_word = 8'h0B;
		16'h9165: out_word = 8'h00;
		16'h9166: out_word = 8'h0A;
		16'h9167: out_word = 8'h00;
		16'h9168: out_word = 8'h09;
		16'h9169: out_word = 8'h00;
		16'h916A: out_word = 8'h09;
		16'h916B: out_word = 8'h00;
		16'h916C: out_word = 8'h08;
		16'h916D: out_word = 8'h00;
		16'h916E: out_word = 8'hDD;
		16'h916F: out_word = 8'h7E;
		16'h9170: out_word = 8'h01;
		16'h9171: out_word = 8'hB7;
		16'h9172: out_word = 8'hF8;
		16'h9173: out_word = 8'hF6;
		16'h9174: out_word = 8'h90;
		16'h9175: out_word = 8'hCD;
		16'h9176: out_word = 8'hA3;
		16'h9177: out_word = 8'h11;
		16'h9178: out_word = 8'hDD;
		16'h9179: out_word = 8'h7E;
		16'h917A: out_word = 8'h00;
		16'h917B: out_word = 8'hCD;
		16'h917C: out_word = 8'hA3;
		16'h917D: out_word = 8'h11;
		16'h917E: out_word = 8'hDD;
		16'h917F: out_word = 8'h7E;
		16'h9180: out_word = 8'h04;
		16'h9181: out_word = 8'hCB;
		16'h9182: out_word = 8'hA7;
		16'h9183: out_word = 8'hCB;
		16'h9184: out_word = 8'h27;
		16'h9185: out_word = 8'hCB;
		16'h9186: out_word = 8'h27;
		16'h9187: out_word = 8'hCB;
		16'h9188: out_word = 8'h27;
		16'h9189: out_word = 8'hCD;
		16'h918A: out_word = 8'hA3;
		16'h918B: out_word = 8'h11;
		16'h918C: out_word = 8'hC9;
		16'h918D: out_word = 8'hDD;
		16'h918E: out_word = 8'h7E;
		16'h918F: out_word = 8'h01;
		16'h9190: out_word = 8'hB7;
		16'h9191: out_word = 8'hF8;
		16'h9192: out_word = 8'hF6;
		16'h9193: out_word = 8'h80;
		16'h9194: out_word = 8'hCD;
		16'h9195: out_word = 8'hA3;
		16'h9196: out_word = 8'h11;
		16'h9197: out_word = 8'hDD;
		16'h9198: out_word = 8'h7E;
		16'h9199: out_word = 8'h00;
		16'h919A: out_word = 8'hCD;
		16'h919B: out_word = 8'hA3;
		16'h919C: out_word = 8'h11;
		16'h919D: out_word = 8'h3E;
		16'h919E: out_word = 8'h40;
		16'h919F: out_word = 8'hCD;
		16'h91A0: out_word = 8'hA3;
		16'h91A1: out_word = 8'h11;
		16'h91A2: out_word = 8'hC9;
		16'h91A3: out_word = 8'h6F;
		16'h91A4: out_word = 8'h01;
		16'h91A5: out_word = 8'hFD;
		16'h91A6: out_word = 8'hFF;
		16'h91A7: out_word = 8'h3E;
		16'h91A8: out_word = 8'h0E;
		16'h91A9: out_word = 8'hED;
		16'h91AA: out_word = 8'h79;
		16'h91AB: out_word = 8'h01;
		16'h91AC: out_word = 8'hFD;
		16'h91AD: out_word = 8'hBF;
		16'h91AE: out_word = 8'h3E;
		16'h91AF: out_word = 8'hFA;
		16'h91B0: out_word = 8'hED;
		16'h91B1: out_word = 8'h79;
		16'h91B2: out_word = 8'h1E;
		16'h91B3: out_word = 8'h03;
		16'h91B4: out_word = 8'h1D;
		16'h91B5: out_word = 8'h20;
		16'h91B6: out_word = 8'hFD;
		16'h91B7: out_word = 8'h00;
		16'h91B8: out_word = 8'h00;
		16'h91B9: out_word = 8'h00;
		16'h91BA: out_word = 8'h00;
		16'h91BB: out_word = 8'h7D;
		16'h91BC: out_word = 8'h16;
		16'h91BD: out_word = 8'h08;
		16'h91BE: out_word = 8'h1F;
		16'h91BF: out_word = 8'h6F;
		16'h91C0: out_word = 8'hD2;
		16'h91C1: out_word = 8'hC9;
		16'h91C2: out_word = 8'h11;
		16'h91C3: out_word = 8'h3E;
		16'h91C4: out_word = 8'hFE;
		16'h91C5: out_word = 8'hED;
		16'h91C6: out_word = 8'h79;
		16'h91C7: out_word = 8'h18;
		16'h91C8: out_word = 8'h06;
		16'h91C9: out_word = 8'h3E;
		16'h91CA: out_word = 8'hFA;
		16'h91CB: out_word = 8'hED;
		16'h91CC: out_word = 8'h79;
		16'h91CD: out_word = 8'h18;
		16'h91CE: out_word = 8'h00;
		16'h91CF: out_word = 8'h1E;
		16'h91D0: out_word = 8'h02;
		16'h91D1: out_word = 8'h1D;
		16'h91D2: out_word = 8'h20;
		16'h91D3: out_word = 8'hFD;
		16'h91D4: out_word = 8'h00;
		16'h91D5: out_word = 8'hC6;
		16'h91D6: out_word = 8'h00;
		16'h91D7: out_word = 8'h7D;
		16'h91D8: out_word = 8'h15;
		16'h91D9: out_word = 8'h20;
		16'h91DA: out_word = 8'hE3;
		16'h91DB: out_word = 8'h00;
		16'h91DC: out_word = 8'h00;
		16'h91DD: out_word = 8'hC6;
		16'h91DE: out_word = 8'h00;
		16'h91DF: out_word = 8'h00;
		16'h91E0: out_word = 8'h00;
		16'h91E1: out_word = 8'h3E;
		16'h91E2: out_word = 8'hFE;
		16'h91E3: out_word = 8'hED;
		16'h91E4: out_word = 8'h79;
		16'h91E5: out_word = 8'h1E;
		16'h91E6: out_word = 8'h06;
		16'h91E7: out_word = 8'h1D;
		16'h91E8: out_word = 8'h20;
		16'h91E9: out_word = 8'hFD;
		16'h91EA: out_word = 8'hC9;
		16'h91EB: out_word = 8'h21;
		16'h91EC: out_word = 8'h66;
		16'h91ED: out_word = 8'h5B;
		16'h91EE: out_word = 8'hCB;
		16'h91EF: out_word = 8'hEE;
		16'h91F0: out_word = 8'h18;
		16'h91F1: out_word = 8'h13;
		16'h91F2: out_word = 8'h21;
		16'h91F3: out_word = 8'h66;
		16'h91F4: out_word = 8'h5B;
		16'h91F5: out_word = 8'hCB;
		16'h91F6: out_word = 8'hE6;
		16'h91F7: out_word = 8'h18;
		16'h91F8: out_word = 8'h0C;
		16'h91F9: out_word = 8'h21;
		16'h91FA: out_word = 8'h66;
		16'h91FB: out_word = 8'h5B;
		16'h91FC: out_word = 8'hCB;
		16'h91FD: out_word = 8'hFE;
		16'h91FE: out_word = 8'h18;
		16'h91FF: out_word = 8'h05;
		16'h9200: out_word = 8'h21;
		16'h9201: out_word = 8'h66;
		16'h9202: out_word = 8'h5B;
		16'h9203: out_word = 8'hCB;
		16'h9204: out_word = 8'hF6;
		16'h9205: out_word = 8'h21;
		16'h9206: out_word = 8'h66;
		16'h9207: out_word = 8'h5B;
		16'h9208: out_word = 8'hCB;
		16'h9209: out_word = 8'h9E;
		16'h920A: out_word = 8'hDF;
		16'h920B: out_word = 8'hFE;
		16'h920C: out_word = 8'h21;
		16'h920D: out_word = 8'hC2;
		16'h920E: out_word = 8'hBE;
		16'h920F: out_word = 8'h13;
		16'h9210: out_word = 8'h21;
		16'h9211: out_word = 8'h66;
		16'h9212: out_word = 8'h5B;
		16'h9213: out_word = 8'hCB;
		16'h9214: out_word = 8'hDE;
		16'h9215: out_word = 8'hE7;
		16'h9216: out_word = 8'hC3;
		16'h9217: out_word = 8'hBE;
		16'h9218: out_word = 8'h13;
		16'h9219: out_word = 8'hCD;
		16'h921A: out_word = 8'hAC;
		16'h921B: out_word = 8'h05;
		16'h921C: out_word = 8'h0B;
		16'h921D: out_word = 8'h22;
		16'h921E: out_word = 8'h74;
		16'h921F: out_word = 8'h5B;
		16'h9220: out_word = 8'hDD;
		16'h9221: out_word = 8'h7E;
		16'h9222: out_word = 8'h00;
		16'h9223: out_word = 8'h32;
		16'h9224: out_word = 8'h71;
		16'h9225: out_word = 8'h5B;
		16'h9226: out_word = 8'hDD;
		16'h9227: out_word = 8'h6E;
		16'h9228: out_word = 8'h0B;
		16'h9229: out_word = 8'hDD;
		16'h922A: out_word = 8'h66;
		16'h922B: out_word = 8'h0C;
		16'h922C: out_word = 8'h22;
		16'h922D: out_word = 8'h72;
		16'h922E: out_word = 8'h5B;
		16'h922F: out_word = 8'hDD;
		16'h9230: out_word = 8'h6E;
		16'h9231: out_word = 8'h0D;
		16'h9232: out_word = 8'hDD;
		16'h9233: out_word = 8'h66;
		16'h9234: out_word = 8'h0E;
		16'h9235: out_word = 8'h22;
		16'h9236: out_word = 8'h78;
		16'h9237: out_word = 8'h5B;
		16'h9238: out_word = 8'hDD;
		16'h9239: out_word = 8'h6E;
		16'h923A: out_word = 8'h0F;
		16'h923B: out_word = 8'hDD;
		16'h923C: out_word = 8'h66;
		16'h923D: out_word = 8'h10;
		16'h923E: out_word = 8'h22;
		16'h923F: out_word = 8'h76;
		16'h9240: out_word = 8'h5B;
		16'h9241: out_word = 8'hB7;
		16'h9242: out_word = 8'h28;
		16'h9243: out_word = 8'h0A;
		16'h9244: out_word = 8'hFE;
		16'h9245: out_word = 8'h03;
		16'h9246: out_word = 8'h28;
		16'h9247: out_word = 8'h06;
		16'h9248: out_word = 8'hDD;
		16'h9249: out_word = 8'h7E;
		16'h924A: out_word = 8'h0E;
		16'h924B: out_word = 8'h32;
		16'h924C: out_word = 8'h76;
		16'h924D: out_word = 8'h5B;
		16'h924E: out_word = 8'hDD;
		16'h924F: out_word = 8'hE5;
		16'h9250: out_word = 8'hE1;
		16'h9251: out_word = 8'h23;
		16'h9252: out_word = 8'h11;
		16'h9253: out_word = 8'h67;
		16'h9254: out_word = 8'h5B;
		16'h9255: out_word = 8'h01;
		16'h9256: out_word = 8'h0A;
		16'h9257: out_word = 8'h00;
		16'h9258: out_word = 8'hED;
		16'h9259: out_word = 8'hB0;
		16'h925A: out_word = 8'h21;
		16'h925B: out_word = 8'h66;
		16'h925C: out_word = 8'h5B;
		16'h925D: out_word = 8'hCB;
		16'h925E: out_word = 8'h6E;
		16'h925F: out_word = 8'hC2;
		16'h9260: out_word = 8'hAD;
		16'h9261: out_word = 8'h1B;
		16'h9262: out_word = 8'h21;
		16'h9263: out_word = 8'h71;
		16'h9264: out_word = 8'h5B;
		16'h9265: out_word = 8'h11;
		16'h9266: out_word = 8'h7A;
		16'h9267: out_word = 8'h5B;
		16'h9268: out_word = 8'h01;
		16'h9269: out_word = 8'h07;
		16'h926A: out_word = 8'h00;
		16'h926B: out_word = 8'hED;
		16'h926C: out_word = 8'hB0;
		16'h926D: out_word = 8'hCD;
		16'h926E: out_word = 8'h2E;
		16'h926F: out_word = 8'h1C;
		16'h9270: out_word = 8'h3A;
		16'h9271: out_word = 8'h7A;
		16'h9272: out_word = 8'h5B;
		16'h9273: out_word = 8'h47;
		16'h9274: out_word = 8'h3A;
		16'h9275: out_word = 8'h71;
		16'h9276: out_word = 8'h5B;
		16'h9277: out_word = 8'hB8;
		16'h9278: out_word = 8'h20;
		16'h9279: out_word = 8'h06;
		16'h927A: out_word = 8'hFE;
		16'h927B: out_word = 8'h03;
		16'h927C: out_word = 8'h28;
		16'h927D: out_word = 8'h12;
		16'h927E: out_word = 8'h38;
		16'h927F: out_word = 8'h04;
		16'h9280: out_word = 8'hCD;
		16'h9281: out_word = 8'hAC;
		16'h9282: out_word = 8'h05;
		16'h9283: out_word = 8'h1D;
		16'h9284: out_word = 8'h3A;
		16'h9285: out_word = 8'h66;
		16'h9286: out_word = 8'h5B;
		16'h9287: out_word = 8'hCB;
		16'h9288: out_word = 8'h77;
		16'h9289: out_word = 8'h20;
		16'h928A: out_word = 8'h3A;
		16'h928B: out_word = 8'hCB;
		16'h928C: out_word = 8'h7F;
		16'h928D: out_word = 8'hCA;
		16'h928E: out_word = 8'hDB;
		16'h928F: out_word = 8'h12;
		16'h9290: out_word = 8'h3A;
		16'h9291: out_word = 8'h66;
		16'h9292: out_word = 8'h5B;
		16'h9293: out_word = 8'hCB;
		16'h9294: out_word = 8'h77;
		16'h9295: out_word = 8'h28;
		16'h9296: out_word = 8'h04;
		16'h9297: out_word = 8'hCD;
		16'h9298: out_word = 8'hAC;
		16'h9299: out_word = 8'h05;
		16'h929A: out_word = 8'h1C;
		16'h929B: out_word = 8'h2A;
		16'h929C: out_word = 8'h7B;
		16'h929D: out_word = 8'h5B;
		16'h929E: out_word = 8'hED;
		16'h929F: out_word = 8'h5B;
		16'h92A0: out_word = 8'h72;
		16'h92A1: out_word = 8'h5B;
		16'h92A2: out_word = 8'h7C;
		16'h92A3: out_word = 8'hB5;
		16'h92A4: out_word = 8'h28;
		16'h92A5: out_word = 8'h08;
		16'h92A6: out_word = 8'hED;
		16'h92A7: out_word = 8'h52;
		16'h92A8: out_word = 8'h30;
		16'h92A9: out_word = 8'h04;
		16'h92AA: out_word = 8'hCD;
		16'h92AB: out_word = 8'hAC;
		16'h92AC: out_word = 8'h05;
		16'h92AD: out_word = 8'h1E;
		16'h92AE: out_word = 8'h2A;
		16'h92AF: out_word = 8'h7D;
		16'h92B0: out_word = 8'h5B;
		16'h92B1: out_word = 8'h7C;
		16'h92B2: out_word = 8'hB5;
		16'h92B3: out_word = 8'h20;
		16'h92B4: out_word = 8'h03;
		16'h92B5: out_word = 8'h2A;
		16'h92B6: out_word = 8'h74;
		16'h92B7: out_word = 8'h5B;
		16'h92B8: out_word = 8'h3A;
		16'h92B9: out_word = 8'h71;
		16'h92BA: out_word = 8'h5B;
		16'h92BB: out_word = 8'hA7;
		16'h92BC: out_word = 8'h20;
		16'h92BD: out_word = 8'h03;
		16'h92BE: out_word = 8'h2A;
		16'h92BF: out_word = 8'h53;
		16'h92C0: out_word = 8'h5C;
		16'h92C1: out_word = 8'hCD;
		16'h92C2: out_word = 8'h7E;
		16'h92C3: out_word = 8'h13;
		16'h92C4: out_word = 8'hC9;
		16'h92C5: out_word = 8'hED;
		16'h92C6: out_word = 8'h4B;
		16'h92C7: out_word = 8'h72;
		16'h92C8: out_word = 8'h5B;
		16'h92C9: out_word = 8'hC5;
		16'h92CA: out_word = 8'h03;
		16'h92CB: out_word = 8'hEF;
		16'h92CC: out_word = 8'h30;
		16'h92CD: out_word = 8'h00;
		16'h92CE: out_word = 8'h36;
		16'h92CF: out_word = 8'h80;
		16'h92D0: out_word = 8'hEB;
		16'h92D1: out_word = 8'hD1;
		16'h92D2: out_word = 8'hE5;
		16'h92D3: out_word = 8'hCD;
		16'h92D4: out_word = 8'h7E;
		16'h92D5: out_word = 8'h13;
		16'h92D6: out_word = 8'hE1;
		16'h92D7: out_word = 8'hEF;
		16'h92D8: out_word = 8'hCE;
		16'h92D9: out_word = 8'h08;
		16'h92DA: out_word = 8'hC9;
		16'h92DB: out_word = 8'hED;
		16'h92DC: out_word = 8'h5B;
		16'h92DD: out_word = 8'h72;
		16'h92DE: out_word = 8'h5B;
		16'h92DF: out_word = 8'h2A;
		16'h92E0: out_word = 8'h7D;
		16'h92E1: out_word = 8'h5B;
		16'h92E2: out_word = 8'hE5;
		16'h92E3: out_word = 8'h7C;
		16'h92E4: out_word = 8'hB5;
		16'h92E5: out_word = 8'h20;
		16'h92E6: out_word = 8'h06;
		16'h92E7: out_word = 8'h13;
		16'h92E8: out_word = 8'h13;
		16'h92E9: out_word = 8'h13;
		16'h92EA: out_word = 8'hEB;
		16'h92EB: out_word = 8'h18;
		16'h92EC: out_word = 8'h09;
		16'h92ED: out_word = 8'h2A;
		16'h92EE: out_word = 8'h7B;
		16'h92EF: out_word = 8'h5B;
		16'h92F0: out_word = 8'hEB;
		16'h92F1: out_word = 8'h37;
		16'h92F2: out_word = 8'hED;
		16'h92F3: out_word = 8'h52;
		16'h92F4: out_word = 8'h38;
		16'h92F5: out_word = 8'h09;
		16'h92F6: out_word = 8'h11;
		16'h92F7: out_word = 8'h05;
		16'h92F8: out_word = 8'h00;
		16'h92F9: out_word = 8'h19;
		16'h92FA: out_word = 8'h44;
		16'h92FB: out_word = 8'h4D;
		16'h92FC: out_word = 8'hEF;
		16'h92FD: out_word = 8'h05;
		16'h92FE: out_word = 8'h1F;
		16'h92FF: out_word = 8'hE1;
		16'h9300: out_word = 8'h3A;
		16'h9301: out_word = 8'h71;
		16'h9302: out_word = 8'h5B;
		16'h9303: out_word = 8'hA7;
		16'h9304: out_word = 8'h28;
		16'h9305: out_word = 8'h2F;
		16'h9306: out_word = 8'h7C;
		16'h9307: out_word = 8'hB5;
		16'h9308: out_word = 8'h28;
		16'h9309: out_word = 8'h0B;
		16'h930A: out_word = 8'h2B;
		16'h930B: out_word = 8'h46;
		16'h930C: out_word = 8'h2B;
		16'h930D: out_word = 8'h4E;
		16'h930E: out_word = 8'h2B;
		16'h930F: out_word = 8'h03;
		16'h9310: out_word = 8'h03;
		16'h9311: out_word = 8'h03;
		16'h9312: out_word = 8'hEF;
		16'h9313: out_word = 8'hE8;
		16'h9314: out_word = 8'h19;
		16'h9315: out_word = 8'h2A;
		16'h9316: out_word = 8'h59;
		16'h9317: out_word = 8'h5C;
		16'h9318: out_word = 8'h2B;
		16'h9319: out_word = 8'hED;
		16'h931A: out_word = 8'h4B;
		16'h931B: out_word = 8'h72;
		16'h931C: out_word = 8'h5B;
		16'h931D: out_word = 8'hC5;
		16'h931E: out_word = 8'h03;
		16'h931F: out_word = 8'h03;
		16'h9320: out_word = 8'h03;
		16'h9321: out_word = 8'h3A;
		16'h9322: out_word = 8'h7F;
		16'h9323: out_word = 8'h5B;
		16'h9324: out_word = 8'hF5;
		16'h9325: out_word = 8'hEF;
		16'h9326: out_word = 8'h55;
		16'h9327: out_word = 8'h16;
		16'h9328: out_word = 8'h23;
		16'h9329: out_word = 8'hF1;
		16'h932A: out_word = 8'h77;
		16'h932B: out_word = 8'hD1;
		16'h932C: out_word = 8'h23;
		16'h932D: out_word = 8'h73;
		16'h932E: out_word = 8'h23;
		16'h932F: out_word = 8'h72;
		16'h9330: out_word = 8'h23;
		16'h9331: out_word = 8'hCD;
		16'h9332: out_word = 8'h7E;
		16'h9333: out_word = 8'h13;
		16'h9334: out_word = 8'hC9;
		16'h9335: out_word = 8'h21;
		16'h9336: out_word = 8'h66;
		16'h9337: out_word = 8'h5B;
		16'h9338: out_word = 8'hCB;
		16'h9339: out_word = 8'h8E;
		16'h933A: out_word = 8'hED;
		16'h933B: out_word = 8'h5B;
		16'h933C: out_word = 8'h53;
		16'h933D: out_word = 8'h5C;
		16'h933E: out_word = 8'h2A;
		16'h933F: out_word = 8'h59;
		16'h9340: out_word = 8'h5C;
		16'h9341: out_word = 8'h2B;
		16'h9342: out_word = 8'hEF;
		16'h9343: out_word = 8'hE5;
		16'h9344: out_word = 8'h19;
		16'h9345: out_word = 8'hED;
		16'h9346: out_word = 8'h4B;
		16'h9347: out_word = 8'h72;
		16'h9348: out_word = 8'h5B;
		16'h9349: out_word = 8'h2A;
		16'h934A: out_word = 8'h53;
		16'h934B: out_word = 8'h5C;
		16'h934C: out_word = 8'hEF;
		16'h934D: out_word = 8'h55;
		16'h934E: out_word = 8'h16;
		16'h934F: out_word = 8'h23;
		16'h9350: out_word = 8'hED;
		16'h9351: out_word = 8'h4B;
		16'h9352: out_word = 8'h76;
		16'h9353: out_word = 8'h5B;
		16'h9354: out_word = 8'h09;
		16'h9355: out_word = 8'h22;
		16'h9356: out_word = 8'h4B;
		16'h9357: out_word = 8'h5C;
		16'h9358: out_word = 8'h3A;
		16'h9359: out_word = 8'h79;
		16'h935A: out_word = 8'h5B;
		16'h935B: out_word = 8'h67;
		16'h935C: out_word = 8'hE6;
		16'h935D: out_word = 8'hC0;
		16'h935E: out_word = 8'h20;
		16'h935F: out_word = 8'h10;
		16'h9360: out_word = 8'h3A;
		16'h9361: out_word = 8'h78;
		16'h9362: out_word = 8'h5B;
		16'h9363: out_word = 8'h6F;
		16'h9364: out_word = 8'h22;
		16'h9365: out_word = 8'h42;
		16'h9366: out_word = 8'h5C;
		16'h9367: out_word = 8'hFD;
		16'h9368: out_word = 8'h36;
		16'h9369: out_word = 8'h0A;
		16'h936A: out_word = 8'h00;
		16'h936B: out_word = 8'h21;
		16'h936C: out_word = 8'h66;
		16'h936D: out_word = 8'h5B;
		16'h936E: out_word = 8'hCB;
		16'h936F: out_word = 8'hCE;
		16'h9370: out_word = 8'h2A;
		16'h9371: out_word = 8'h53;
		16'h9372: out_word = 8'h5C;
		16'h9373: out_word = 8'hED;
		16'h9374: out_word = 8'h5B;
		16'h9375: out_word = 8'h72;
		16'h9376: out_word = 8'h5B;
		16'h9377: out_word = 8'h2B;
		16'h9378: out_word = 8'h22;
		16'h9379: out_word = 8'h57;
		16'h937A: out_word = 8'h5C;
		16'h937B: out_word = 8'h23;
		16'h937C: out_word = 8'h18;
		16'h937D: out_word = 8'hB3;
		16'h937E: out_word = 8'h7A;
		16'h937F: out_word = 8'hB3;
		16'h9380: out_word = 8'hC8;
		16'h9381: out_word = 8'hCD;
		16'h9382: out_word = 8'h4B;
		16'h9383: out_word = 8'h1C;
		16'h9384: out_word = 8'hC9;
		16'h9385: out_word = 8'hEF;
		16'h9386: out_word = 8'h8C;
		16'h9387: out_word = 8'h1C;
		16'h9388: out_word = 8'hFD;
		16'h9389: out_word = 8'hCB;
		16'h938A: out_word = 8'h01;
		16'h938B: out_word = 8'h7E;
		16'h938C: out_word = 8'hC8;
		16'h938D: out_word = 8'hF5;
		16'h938E: out_word = 8'hEF;
		16'h938F: out_word = 8'hF1;
		16'h9390: out_word = 8'h2B;
		16'h9391: out_word = 8'hF1;
		16'h9392: out_word = 8'hC9;
		16'h9393: out_word = 8'hE7;
		16'h9394: out_word = 8'hCD;
		16'h9395: out_word = 8'h85;
		16'h9396: out_word = 8'h13;
		16'h9397: out_word = 8'hC8;
		16'h9398: out_word = 8'hF5;
		16'h9399: out_word = 8'h79;
		16'h939A: out_word = 8'hB0;
		16'h939B: out_word = 8'h28;
		16'h939C: out_word = 8'h1D;
		16'h939D: out_word = 8'h21;
		16'h939E: out_word = 8'h0A;
		16'h939F: out_word = 8'h00;
		16'h93A0: out_word = 8'hED;
		16'h93A1: out_word = 8'h42;
		16'h93A2: out_word = 8'h38;
		16'h93A3: out_word = 8'h16;
		16'h93A4: out_word = 8'hD5;
		16'h93A5: out_word = 8'hC5;
		16'h93A6: out_word = 8'h21;
		16'h93A7: out_word = 8'h67;
		16'h93A8: out_word = 8'h5B;
		16'h93A9: out_word = 8'h06;
		16'h93AA: out_word = 8'h0A;
		16'h93AB: out_word = 8'h3E;
		16'h93AC: out_word = 8'h20;
		16'h93AD: out_word = 8'h77;
		16'h93AE: out_word = 8'h23;
		16'h93AF: out_word = 8'h10;
		16'h93B0: out_word = 8'hFC;
		16'h93B1: out_word = 8'hC1;
		16'h93B2: out_word = 8'hE1;
		16'h93B3: out_word = 8'h11;
		16'h93B4: out_word = 8'h67;
		16'h93B5: out_word = 8'h5B;
		16'h93B6: out_word = 8'hED;
		16'h93B7: out_word = 8'hB0;
		16'h93B8: out_word = 8'hF1;
		16'h93B9: out_word = 8'hC9;
		16'h93BA: out_word = 8'hCD;
		16'h93BB: out_word = 8'hAC;
		16'h93BC: out_word = 8'h05;
		16'h93BD: out_word = 8'h21;
		16'h93BE: out_word = 8'hEF;
		16'h93BF: out_word = 8'h8C;
		16'h93C0: out_word = 8'h1C;
		16'h93C1: out_word = 8'hFD;
		16'h93C2: out_word = 8'hCB;
		16'h93C3: out_word = 8'h01;
		16'h93C4: out_word = 8'h7E;
		16'h93C5: out_word = 8'h28;
		16'h93C6: out_word = 8'h40;
		16'h93C7: out_word = 8'h01;
		16'h93C8: out_word = 8'h11;
		16'h93C9: out_word = 8'h00;
		16'h93CA: out_word = 8'h3A;
		16'h93CB: out_word = 8'h74;
		16'h93CC: out_word = 8'h5C;
		16'h93CD: out_word = 8'hA7;
		16'h93CE: out_word = 8'h28;
		16'h93CF: out_word = 8'h02;
		16'h93D0: out_word = 8'h0E;
		16'h93D1: out_word = 8'h22;
		16'h93D2: out_word = 8'hEF;
		16'h93D3: out_word = 8'h30;
		16'h93D4: out_word = 8'h00;
		16'h93D5: out_word = 8'hD5;
		16'h93D6: out_word = 8'hDD;
		16'h93D7: out_word = 8'hE1;
		16'h93D8: out_word = 8'h06;
		16'h93D9: out_word = 8'h0B;
		16'h93DA: out_word = 8'h3E;
		16'h93DB: out_word = 8'h20;
		16'h93DC: out_word = 8'h12;
		16'h93DD: out_word = 8'h13;
		16'h93DE: out_word = 8'h10;
		16'h93DF: out_word = 8'hFC;
		16'h93E0: out_word = 8'hDD;
		16'h93E1: out_word = 8'h36;
		16'h93E2: out_word = 8'h01;
		16'h93E3: out_word = 8'hFF;
		16'h93E4: out_word = 8'hEF;
		16'h93E5: out_word = 8'hF1;
		16'h93E6: out_word = 8'h2B;
		16'h93E7: out_word = 8'h21;
		16'h93E8: out_word = 8'hF6;
		16'h93E9: out_word = 8'hFF;
		16'h93EA: out_word = 8'h0B;
		16'h93EB: out_word = 8'h09;
		16'h93EC: out_word = 8'h03;
		16'h93ED: out_word = 8'h30;
		16'h93EE: out_word = 8'h11;
		16'h93EF: out_word = 8'h3A;
		16'h93F0: out_word = 8'h74;
		16'h93F1: out_word = 8'h5C;
		16'h93F2: out_word = 8'hA7;
		16'h93F3: out_word = 8'h20;
		16'h93F4: out_word = 8'h04;
		16'h93F5: out_word = 8'hCD;
		16'h93F6: out_word = 8'hAC;
		16'h93F7: out_word = 8'h05;
		16'h93F8: out_word = 8'h0E;
		16'h93F9: out_word = 8'h78;
		16'h93FA: out_word = 8'hB1;
		16'h93FB: out_word = 8'h28;
		16'h93FC: out_word = 8'h0A;
		16'h93FD: out_word = 8'h01;
		16'h93FE: out_word = 8'h0A;
		16'h93FF: out_word = 8'h00;
		16'h9400: out_word = 8'hDD;
		16'h9401: out_word = 8'hE5;
		16'h9402: out_word = 8'hE1;
		16'h9403: out_word = 8'h23;
		16'h9404: out_word = 8'hEB;
		16'h9405: out_word = 8'hED;
		16'h9406: out_word = 8'hB0;
		16'h9407: out_word = 8'hDF;
		16'h9408: out_word = 8'hFE;
		16'h9409: out_word = 8'hE4;
		16'h940A: out_word = 8'h20;
		16'h940B: out_word = 8'h53;
		16'h940C: out_word = 8'h3A;
		16'h940D: out_word = 8'h74;
		16'h940E: out_word = 8'h5C;
		16'h940F: out_word = 8'hFE;
		16'h9410: out_word = 8'h03;
		16'h9411: out_word = 8'hCA;
		16'h9412: out_word = 8'h19;
		16'h9413: out_word = 8'h12;
		16'h9414: out_word = 8'hE7;
		16'h9415: out_word = 8'hEF;
		16'h9416: out_word = 8'hB2;
		16'h9417: out_word = 8'h28;
		16'h9418: out_word = 8'h30;
		16'h9419: out_word = 8'h15;
		16'h941A: out_word = 8'h21;
		16'h941B: out_word = 8'h00;
		16'h941C: out_word = 8'h00;
		16'h941D: out_word = 8'hFD;
		16'h941E: out_word = 8'hCB;
		16'h941F: out_word = 8'h01;
		16'h9420: out_word = 8'h76;
		16'h9421: out_word = 8'h28;
		16'h9422: out_word = 8'h02;
		16'h9423: out_word = 8'hCB;
		16'h9424: out_word = 8'hF9;
		16'h9425: out_word = 8'h3A;
		16'h9426: out_word = 8'h74;
		16'h9427: out_word = 8'h5C;
		16'h9428: out_word = 8'h3D;
		16'h9429: out_word = 8'h28;
		16'h942A: out_word = 8'h19;
		16'h942B: out_word = 8'hCD;
		16'h942C: out_word = 8'hAC;
		16'h942D: out_word = 8'h05;
		16'h942E: out_word = 8'h01;
		16'h942F: out_word = 8'hC2;
		16'h9430: out_word = 8'h19;
		16'h9431: out_word = 8'h12;
		16'h9432: out_word = 8'hFD;
		16'h9433: out_word = 8'hCB;
		16'h9434: out_word = 8'h01;
		16'h9435: out_word = 8'h7E;
		16'h9436: out_word = 8'h28;
		16'h9437: out_word = 8'h19;
		16'h9438: out_word = 8'h4E;
		16'h9439: out_word = 8'h23;
		16'h943A: out_word = 8'h7E;
		16'h943B: out_word = 8'hDD;
		16'h943C: out_word = 8'h77;
		16'h943D: out_word = 8'h0B;
		16'h943E: out_word = 8'h23;
		16'h943F: out_word = 8'h7E;
		16'h9440: out_word = 8'hDD;
		16'h9441: out_word = 8'h77;
		16'h9442: out_word = 8'h0C;
		16'h9443: out_word = 8'h23;
		16'h9444: out_word = 8'hDD;
		16'h9445: out_word = 8'h71;
		16'h9446: out_word = 8'h0E;
		16'h9447: out_word = 8'h3E;
		16'h9448: out_word = 8'h01;
		16'h9449: out_word = 8'hCB;
		16'h944A: out_word = 8'h71;
		16'h944B: out_word = 8'h28;
		16'h944C: out_word = 8'h01;
		16'h944D: out_word = 8'h3C;
		16'h944E: out_word = 8'hDD;
		16'h944F: out_word = 8'h77;
		16'h9450: out_word = 8'h00;
		16'h9451: out_word = 8'hEB;
		16'h9452: out_word = 8'hE7;
		16'h9453: out_word = 8'hFE;
		16'h9454: out_word = 8'h29;
		16'h9455: out_word = 8'h20;
		16'h9456: out_word = 8'hD8;
		16'h9457: out_word = 8'hE7;
		16'h9458: out_word = 8'hCD;
		16'h9459: out_word = 8'hA1;
		16'h945A: out_word = 8'h18;
		16'h945B: out_word = 8'hEB;
		16'h945C: out_word = 8'hC3;
		16'h945D: out_word = 8'h19;
		16'h945E: out_word = 8'h15;
		16'h945F: out_word = 8'hFE;
		16'h9460: out_word = 8'hAA;
		16'h9461: out_word = 8'h20;
		16'h9462: out_word = 8'h1F;
		16'h9463: out_word = 8'h3A;
		16'h9464: out_word = 8'h74;
		16'h9465: out_word = 8'h5C;
		16'h9466: out_word = 8'hFE;
		16'h9467: out_word = 8'h03;
		16'h9468: out_word = 8'hCA;
		16'h9469: out_word = 8'h19;
		16'h946A: out_word = 8'h12;
		16'h946B: out_word = 8'hE7;
		16'h946C: out_word = 8'hCD;
		16'h946D: out_word = 8'hA1;
		16'h946E: out_word = 8'h18;
		16'h946F: out_word = 8'hDD;
		16'h9470: out_word = 8'h36;
		16'h9471: out_word = 8'h0B;
		16'h9472: out_word = 8'h00;
		16'h9473: out_word = 8'hDD;
		16'h9474: out_word = 8'h36;
		16'h9475: out_word = 8'h0C;
		16'h9476: out_word = 8'h1B;
		16'h9477: out_word = 8'h21;
		16'h9478: out_word = 8'h00;
		16'h9479: out_word = 8'h40;
		16'h947A: out_word = 8'hDD;
		16'h947B: out_word = 8'h75;
		16'h947C: out_word = 8'h0D;
		16'h947D: out_word = 8'hDD;
		16'h947E: out_word = 8'h74;
		16'h947F: out_word = 8'h0E;
		16'h9480: out_word = 8'h18;
		16'h9481: out_word = 8'h4D;
		16'h9482: out_word = 8'hFE;
		16'h9483: out_word = 8'hAF;
		16'h9484: out_word = 8'h20;
		16'h9485: out_word = 8'h4F;
		16'h9486: out_word = 8'h3A;
		16'h9487: out_word = 8'h74;
		16'h9488: out_word = 8'h5C;
		16'h9489: out_word = 8'hFE;
		16'h948A: out_word = 8'h03;
		16'h948B: out_word = 8'hCA;
		16'h948C: out_word = 8'h19;
		16'h948D: out_word = 8'h12;
		16'h948E: out_word = 8'hE7;
		16'h948F: out_word = 8'hEF;
		16'h9490: out_word = 8'h48;
		16'h9491: out_word = 8'h20;
		16'h9492: out_word = 8'h20;
		16'h9493: out_word = 8'h0C;
		16'h9494: out_word = 8'h3A;
		16'h9495: out_word = 8'h74;
		16'h9496: out_word = 8'h5C;
		16'h9497: out_word = 8'hA7;
		16'h9498: out_word = 8'hCA;
		16'h9499: out_word = 8'h19;
		16'h949A: out_word = 8'h12;
		16'h949B: out_word = 8'hEF;
		16'h949C: out_word = 8'hE6;
		16'h949D: out_word = 8'h1C;
		16'h949E: out_word = 8'h18;
		16'h949F: out_word = 8'h0F;
		16'h94A0: out_word = 8'hEF;
		16'h94A1: out_word = 8'h82;
		16'h94A2: out_word = 8'h1C;
		16'h94A3: out_word = 8'hDF;
		16'h94A4: out_word = 8'hFE;
		16'h94A5: out_word = 8'h2C;
		16'h94A6: out_word = 8'h28;
		16'h94A7: out_word = 8'h0C;
		16'h94A8: out_word = 8'h3A;
		16'h94A9: out_word = 8'h74;
		16'h94AA: out_word = 8'h5C;
		16'h94AB: out_word = 8'hA7;
		16'h94AC: out_word = 8'hCA;
		16'h94AD: out_word = 8'h19;
		16'h94AE: out_word = 8'h12;
		16'h94AF: out_word = 8'hEF;
		16'h94B0: out_word = 8'hE6;
		16'h94B1: out_word = 8'h1C;
		16'h94B2: out_word = 8'h18;
		16'h94B3: out_word = 8'h04;
		16'h94B4: out_word = 8'hE7;
		16'h94B5: out_word = 8'hEF;
		16'h94B6: out_word = 8'h82;
		16'h94B7: out_word = 8'h1C;
		16'h94B8: out_word = 8'hCD;
		16'h94B9: out_word = 8'hA1;
		16'h94BA: out_word = 8'h18;
		16'h94BB: out_word = 8'hEF;
		16'h94BC: out_word = 8'h99;
		16'h94BD: out_word = 8'h1E;
		16'h94BE: out_word = 8'hDD;
		16'h94BF: out_word = 8'h71;
		16'h94C0: out_word = 8'h0B;
		16'h94C1: out_word = 8'hDD;
		16'h94C2: out_word = 8'h70;
		16'h94C3: out_word = 8'h0C;
		16'h94C4: out_word = 8'hEF;
		16'h94C5: out_word = 8'h99;
		16'h94C6: out_word = 8'h1E;
		16'h94C7: out_word = 8'hDD;
		16'h94C8: out_word = 8'h71;
		16'h94C9: out_word = 8'h0D;
		16'h94CA: out_word = 8'hDD;
		16'h94CB: out_word = 8'h70;
		16'h94CC: out_word = 8'h0E;
		16'h94CD: out_word = 8'h60;
		16'h94CE: out_word = 8'h69;
		16'h94CF: out_word = 8'hDD;
		16'h94D0: out_word = 8'h36;
		16'h94D1: out_word = 8'h00;
		16'h94D2: out_word = 8'h03;
		16'h94D3: out_word = 8'h18;
		16'h94D4: out_word = 8'h44;
		16'h94D5: out_word = 8'hFE;
		16'h94D6: out_word = 8'hCA;
		16'h94D7: out_word = 8'h28;
		16'h94D8: out_word = 8'h09;
		16'h94D9: out_word = 8'hCD;
		16'h94DA: out_word = 8'hA1;
		16'h94DB: out_word = 8'h18;
		16'h94DC: out_word = 8'hDD;
		16'h94DD: out_word = 8'h36;
		16'h94DE: out_word = 8'h0E;
		16'h94DF: out_word = 8'h80;
		16'h94E0: out_word = 8'h18;
		16'h94E1: out_word = 8'h17;
		16'h94E2: out_word = 8'h3A;
		16'h94E3: out_word = 8'h74;
		16'h94E4: out_word = 8'h5C;
		16'h94E5: out_word = 8'hA7;
		16'h94E6: out_word = 8'hC2;
		16'h94E7: out_word = 8'h19;
		16'h94E8: out_word = 8'h12;
		16'h94E9: out_word = 8'hE7;
		16'h94EA: out_word = 8'hEF;
		16'h94EB: out_word = 8'h82;
		16'h94EC: out_word = 8'h1C;
		16'h94ED: out_word = 8'hCD;
		16'h94EE: out_word = 8'hA1;
		16'h94EF: out_word = 8'h18;
		16'h94F0: out_word = 8'hEF;
		16'h94F1: out_word = 8'h99;
		16'h94F2: out_word = 8'h1E;
		16'h94F3: out_word = 8'hDD;
		16'h94F4: out_word = 8'h71;
		16'h94F5: out_word = 8'h0D;
		16'h94F6: out_word = 8'hDD;
		16'h94F7: out_word = 8'h70;
		16'h94F8: out_word = 8'h0E;
		16'h94F9: out_word = 8'hDD;
		16'h94FA: out_word = 8'h36;
		16'h94FB: out_word = 8'h00;
		16'h94FC: out_word = 8'h00;
		16'h94FD: out_word = 8'h2A;
		16'h94FE: out_word = 8'h59;
		16'h94FF: out_word = 8'h5C;
		16'h9500: out_word = 8'hED;
		16'h9501: out_word = 8'h5B;
		16'h9502: out_word = 8'h53;
		16'h9503: out_word = 8'h5C;
		16'h9504: out_word = 8'h37;
		16'h9505: out_word = 8'hED;
		16'h9506: out_word = 8'h52;
		16'h9507: out_word = 8'hDD;
		16'h9508: out_word = 8'h75;
		16'h9509: out_word = 8'h0B;
		16'h950A: out_word = 8'hDD;
		16'h950B: out_word = 8'h74;
		16'h950C: out_word = 8'h0C;
		16'h950D: out_word = 8'h2A;
		16'h950E: out_word = 8'h4B;
		16'h950F: out_word = 8'h5C;
		16'h9510: out_word = 8'hED;
		16'h9511: out_word = 8'h52;
		16'h9512: out_word = 8'hDD;
		16'h9513: out_word = 8'h75;
		16'h9514: out_word = 8'h0F;
		16'h9515: out_word = 8'hDD;
		16'h9516: out_word = 8'h74;
		16'h9517: out_word = 8'h10;
		16'h9518: out_word = 8'hEB;
		16'h9519: out_word = 8'h3A;
		16'h951A: out_word = 8'h66;
		16'h951B: out_word = 8'h5B;
		16'h951C: out_word = 8'hCB;
		16'h951D: out_word = 8'h5F;
		16'h951E: out_word = 8'hC2;
		16'h951F: out_word = 8'h1D;
		16'h9520: out_word = 8'h12;
		16'h9521: out_word = 8'h3A;
		16'h9522: out_word = 8'h74;
		16'h9523: out_word = 8'h5C;
		16'h9524: out_word = 8'hA7;
		16'h9525: out_word = 8'h20;
		16'h9526: out_word = 8'h04;
		16'h9527: out_word = 8'hEF;
		16'h9528: out_word = 8'h70;
		16'h9529: out_word = 8'h09;
		16'h952A: out_word = 8'hC9;
		16'h952B: out_word = 8'hEF;
		16'h952C: out_word = 8'h61;
		16'h952D: out_word = 8'h07;
		16'h952E: out_word = 8'hC9;
		16'h952F: out_word = 8'h21;
		16'h9530: out_word = 8'hF5;
		16'h9531: out_word = 8'hEE;
		16'h9532: out_word = 8'hCB;
		16'h9533: out_word = 8'h86;
		16'h9534: out_word = 8'hCB;
		16'h9535: out_word = 8'hCE;
		16'h9536: out_word = 8'h2A;
		16'h9537: out_word = 8'h49;
		16'h9538: out_word = 8'h5C;
		16'h9539: out_word = 8'h7C;
		16'h953A: out_word = 8'hB5;
		16'h953B: out_word = 8'h20;
		16'h953C: out_word = 8'h03;
		16'h953D: out_word = 8'h22;
		16'h953E: out_word = 8'h06;
		16'h953F: out_word = 8'hEC;
		16'h9540: out_word = 8'h3A;
		16'h9541: out_word = 8'hDB;
		16'h9542: out_word = 8'hF9;
		16'h9543: out_word = 8'hF5;
		16'h9544: out_word = 8'h2A;
		16'h9545: out_word = 8'h9A;
		16'h9546: out_word = 8'hFC;
		16'h9547: out_word = 8'hCD;
		16'h9548: out_word = 8'h4A;
		16'h9549: out_word = 8'h33;
		16'h954A: out_word = 8'h22;
		16'h954B: out_word = 8'hD7;
		16'h954C: out_word = 8'hF9;
		16'h954D: out_word = 8'hCD;
		16'h954E: out_word = 8'h22;
		16'h954F: out_word = 8'h32;
		16'h9550: out_word = 8'hCD;
		16'h9551: out_word = 8'hD6;
		16'h9552: out_word = 8'h30;
		16'h9553: out_word = 8'hF1;
		16'h9554: out_word = 8'hB7;
		16'h9555: out_word = 8'h28;
		16'h9556: out_word = 8'h0C;
		16'h9557: out_word = 8'hF5;
		16'h9558: out_word = 8'hCD;
		16'h9559: out_word = 8'hDF;
		16'h955A: out_word = 8'h30;
		16'h955B: out_word = 8'hEB;
		16'h955C: out_word = 8'hCD;
		16'h955D: out_word = 8'h6A;
		16'h955E: out_word = 8'h32;
		16'h955F: out_word = 8'hF1;
		16'h9560: out_word = 8'h3D;
		16'h9561: out_word = 8'h18;
		16'h9562: out_word = 8'hF1;
		16'h9563: out_word = 8'h0E;
		16'h9564: out_word = 8'h00;
		16'h9565: out_word = 8'hCD;
		16'h9566: out_word = 8'hB4;
		16'h9567: out_word = 8'h30;
		16'h9568: out_word = 8'h41;
		16'h9569: out_word = 8'h3A;
		16'h956A: out_word = 8'h15;
		16'h956B: out_word = 8'hEC;
		16'h956C: out_word = 8'h4F;
		16'h956D: out_word = 8'hC5;
		16'h956E: out_word = 8'hD5;
		16'h956F: out_word = 8'hCD;
		16'h9570: out_word = 8'hDF;
		16'h9571: out_word = 8'h30;
		16'h9572: out_word = 8'h3A;
		16'h9573: out_word = 8'hF5;
		16'h9574: out_word = 8'hEE;
		16'h9575: out_word = 8'hCB;
		16'h9576: out_word = 8'h4F;
		16'h9577: out_word = 8'h28;
		16'h9578: out_word = 8'h1D;
		16'h9579: out_word = 8'hD5;
		16'h957A: out_word = 8'hE5;
		16'h957B: out_word = 8'h11;
		16'h957C: out_word = 8'h20;
		16'h957D: out_word = 8'h00;
		16'h957E: out_word = 8'h19;
		16'h957F: out_word = 8'hCB;
		16'h9580: out_word = 8'h46;
		16'h9581: out_word = 8'h28;
		16'h9582: out_word = 8'h11;
		16'h9583: out_word = 8'h23;
		16'h9584: out_word = 8'h56;
		16'h9585: out_word = 8'h23;
		16'h9586: out_word = 8'h5E;
		16'h9587: out_word = 8'hB7;
		16'h9588: out_word = 8'h2A;
		16'h9589: out_word = 8'h49;
		16'h958A: out_word = 8'h5C;
		16'h958B: out_word = 8'hED;
		16'h958C: out_word = 8'h52;
		16'h958D: out_word = 8'h20;
		16'h958E: out_word = 8'h05;
		16'h958F: out_word = 8'h21;
		16'h9590: out_word = 8'hF5;
		16'h9591: out_word = 8'hEE;
		16'h9592: out_word = 8'hCB;
		16'h9593: out_word = 8'hC6;
		16'h9594: out_word = 8'hE1;
		16'h9595: out_word = 8'hD1;
		16'h9596: out_word = 8'hC5;
		16'h9597: out_word = 8'hE5;
		16'h9598: out_word = 8'h01;
		16'h9599: out_word = 8'h23;
		16'h959A: out_word = 8'h00;
		16'h959B: out_word = 8'hED;
		16'h959C: out_word = 8'hB0;
		16'h959D: out_word = 8'hE1;
		16'h959E: out_word = 8'hC1;
		16'h959F: out_word = 8'hD5;
		16'h95A0: out_word = 8'hC5;
		16'h95A1: out_word = 8'hEB;
		16'h95A2: out_word = 8'h21;
		16'h95A3: out_word = 8'hF5;
		16'h95A4: out_word = 8'hEE;
		16'h95A5: out_word = 8'hCB;
		16'h95A6: out_word = 8'h46;
		16'h95A7: out_word = 8'h28;
		16'h95A8: out_word = 8'h2A;
		16'h95A9: out_word = 8'h06;
		16'h95AA: out_word = 8'h00;
		16'h95AB: out_word = 8'h2A;
		16'h95AC: out_word = 8'h06;
		16'h95AD: out_word = 8'hEC;
		16'h95AE: out_word = 8'h7C;
		16'h95AF: out_word = 8'hB5;
		16'h95B0: out_word = 8'h28;
		16'h95B1: out_word = 8'h0E;
		16'h95B2: out_word = 8'hE5;
		16'h95B3: out_word = 8'hCD;
		16'h95B4: out_word = 8'h41;
		16'h95B5: out_word = 8'h2E;
		16'h95B6: out_word = 8'hE1;
		16'h95B7: out_word = 8'h30;
		16'h95B8: out_word = 8'h12;
		16'h95B9: out_word = 8'h2B;
		16'h95BA: out_word = 8'h04;
		16'h95BB: out_word = 8'h22;
		16'h95BC: out_word = 8'h06;
		16'h95BD: out_word = 8'hEC;
		16'h95BE: out_word = 8'h18;
		16'h95BF: out_word = 8'hEB;
		16'h95C0: out_word = 8'hCD;
		16'h95C1: out_word = 8'h41;
		16'h95C2: out_word = 8'h2E;
		16'h95C3: out_word = 8'hD4;
		16'h95C4: out_word = 8'h63;
		16'h95C5: out_word = 8'h2E;
		16'h95C6: out_word = 8'h21;
		16'h95C7: out_word = 8'hF5;
		16'h95C8: out_word = 8'hEE;
		16'h95C9: out_word = 8'h36;
		16'h95CA: out_word = 8'h00;
		16'h95CB: out_word = 8'h78;
		16'h95CC: out_word = 8'hC1;
		16'h95CD: out_word = 8'hC5;
		16'h95CE: out_word = 8'h48;
		16'h95CF: out_word = 8'h47;
		16'h95D0: out_word = 8'hCD;
		16'h95D1: out_word = 8'h11;
		16'h95D2: out_word = 8'h2A;
		16'h95D3: out_word = 8'hC1;
		16'h95D4: out_word = 8'hD1;
		16'h95D5: out_word = 8'h79;
		16'h95D6: out_word = 8'h04;
		16'h95D7: out_word = 8'hB8;
		16'h95D8: out_word = 8'h30;
		16'h95D9: out_word = 8'h95;
		16'h95DA: out_word = 8'h3A;
		16'h95DB: out_word = 8'hF5;
		16'h95DC: out_word = 8'hEE;
		16'h95DD: out_word = 8'hCB;
		16'h95DE: out_word = 8'h4F;
		16'h95DF: out_word = 8'h28;
		16'h95E0: out_word = 8'h21;
		16'h95E1: out_word = 8'hCB;
		16'h95E2: out_word = 8'h47;
		16'h95E3: out_word = 8'h20;
		16'h95E4: out_word = 8'h1D;
		16'h95E5: out_word = 8'h2A;
		16'h95E6: out_word = 8'h49;
		16'h95E7: out_word = 8'h5C;
		16'h95E8: out_word = 8'h7C;
		16'h95E9: out_word = 8'hB5;
		16'h95EA: out_word = 8'h28;
		16'h95EB: out_word = 8'h08;
		16'h95EC: out_word = 8'h22;
		16'h95ED: out_word = 8'h9A;
		16'h95EE: out_word = 8'hFC;
		16'h95EF: out_word = 8'hCD;
		16'h95F0: out_word = 8'h22;
		16'h95F1: out_word = 8'h32;
		16'h95F2: out_word = 8'h18;
		16'h95F3: out_word = 8'h09;
		16'h95F4: out_word = 8'h22;
		16'h95F5: out_word = 8'h9A;
		16'h95F6: out_word = 8'hFC;
		16'h95F7: out_word = 8'hCD;
		16'h95F8: out_word = 8'h52;
		16'h95F9: out_word = 8'h33;
		16'h95FA: out_word = 8'h22;
		16'h95FB: out_word = 8'h49;
		16'h95FC: out_word = 8'h5C;
		16'h95FD: out_word = 8'hD1;
		16'h95FE: out_word = 8'hC1;
		16'h95FF: out_word = 8'hC3;
		16'h9600: out_word = 8'h36;
		16'h9601: out_word = 8'h15;
		16'h9602: out_word = 8'hD1;
		16'h9603: out_word = 8'hC1;
		16'h9604: out_word = 8'hBF;
		16'h9605: out_word = 8'hF5;
		16'h9606: out_word = 8'h79;
		16'h9607: out_word = 8'h48;
		16'h9608: out_word = 8'hCD;
		16'h9609: out_word = 8'hB4;
		16'h960A: out_word = 8'h30;
		16'h960B: out_word = 8'hEB;
		16'h960C: out_word = 8'hF5;
		16'h960D: out_word = 8'hCD;
		16'h960E: out_word = 8'h04;
		16'h960F: out_word = 8'h36;
		16'h9610: out_word = 8'hF1;
		16'h9611: out_word = 8'h11;
		16'h9612: out_word = 8'h23;
		16'h9613: out_word = 8'h00;
		16'h9614: out_word = 8'h19;
		16'h9615: out_word = 8'h0C;
		16'h9616: out_word = 8'hB9;
		16'h9617: out_word = 8'h30;
		16'h9618: out_word = 8'hF3;
		16'h9619: out_word = 8'hF1;
		16'h961A: out_word = 8'hC8;
		16'h961B: out_word = 8'hCD;
		16'h961C: out_word = 8'h07;
		16'h961D: out_word = 8'h2A;
		16'h961E: out_word = 8'hCD;
		16'h961F: out_word = 8'h78;
		16'h9620: out_word = 8'h2B;
		16'h9621: out_word = 8'h2A;
		16'h9622: out_word = 8'h06;
		16'h9623: out_word = 8'hEC;
		16'h9624: out_word = 8'h2B;
		16'h9625: out_word = 8'h7C;
		16'h9626: out_word = 8'hB5;
		16'h9627: out_word = 8'h22;
		16'h9628: out_word = 8'h06;
		16'h9629: out_word = 8'hEC;
		16'h962A: out_word = 8'h20;
		16'h962B: out_word = 8'hF2;
		16'h962C: out_word = 8'hC3;
		16'h962D: out_word = 8'h11;
		16'h962E: out_word = 8'h2A;
		16'h962F: out_word = 8'hC9;
		16'h9630: out_word = 8'h06;
		16'h9631: out_word = 8'h00;
		16'h9632: out_word = 8'h3A;
		16'h9633: out_word = 8'h15;
		16'h9634: out_word = 8'hEC;
		16'h9635: out_word = 8'h57;
		16'h9636: out_word = 8'hC3;
		16'h9637: out_word = 8'h5E;
		16'h9638: out_word = 8'h3B;
		16'h9639: out_word = 8'h06;
		16'h963A: out_word = 8'h00;
		16'h963B: out_word = 8'hE5;
		16'h963C: out_word = 8'h48;
		16'h963D: out_word = 8'hCD;
		16'h963E: out_word = 8'hB4;
		16'h963F: out_word = 8'h30;
		16'h9640: out_word = 8'hCD;
		16'h9641: out_word = 8'h6A;
		16'h9642: out_word = 8'h32;
		16'h9643: out_word = 8'hE1;
		16'h9644: out_word = 8'hD0;
		16'h9645: out_word = 8'hCD;
		16'h9646: out_word = 8'hDF;
		16'h9647: out_word = 8'h30;
		16'h9648: out_word = 8'hC5;
		16'h9649: out_word = 8'hE5;
		16'h964A: out_word = 8'h21;
		16'h964B: out_word = 8'h23;
		16'h964C: out_word = 8'h00;
		16'h964D: out_word = 8'h19;
		16'h964E: out_word = 8'h3A;
		16'h964F: out_word = 8'h15;
		16'h9650: out_word = 8'hEC;
		16'h9651: out_word = 8'h4F;
		16'h9652: out_word = 8'hB8;
		16'h9653: out_word = 8'h28;
		16'h9654: out_word = 8'h0E;
		16'h9655: out_word = 8'hC5;
		16'h9656: out_word = 8'hC5;
		16'h9657: out_word = 8'h01;
		16'h9658: out_word = 8'h23;
		16'h9659: out_word = 8'h00;
		16'h965A: out_word = 8'hED;
		16'h965B: out_word = 8'hB0;
		16'h965C: out_word = 8'hC1;
		16'h965D: out_word = 8'h79;
		16'h965E: out_word = 8'h04;
		16'h965F: out_word = 8'hB8;
		16'h9660: out_word = 8'h20;
		16'h9661: out_word = 8'hF4;
		16'h9662: out_word = 8'hC1;
		16'h9663: out_word = 8'hE1;
		16'h9664: out_word = 8'hCD;
		16'h9665: out_word = 8'h18;
		16'h9666: out_word = 8'h36;
		16'h9667: out_word = 8'h01;
		16'h9668: out_word = 8'h23;
		16'h9669: out_word = 8'h00;
		16'h966A: out_word = 8'hED;
		16'h966B: out_word = 8'hB0;
		16'h966C: out_word = 8'h37;
		16'h966D: out_word = 8'hC1;
		16'h966E: out_word = 8'hC9;
		16'h966F: out_word = 8'h06;
		16'h9670: out_word = 8'h00;
		16'h9671: out_word = 8'hCD;
		16'h9672: out_word = 8'h2B;
		16'h9673: out_word = 8'h32;
		16'h9674: out_word = 8'hD0;
		16'h9675: out_word = 8'hC5;
		16'h9676: out_word = 8'hE5;
		16'h9677: out_word = 8'h3A;
		16'h9678: out_word = 8'h15;
		16'h9679: out_word = 8'hEC;
		16'h967A: out_word = 8'h4F;
		16'h967B: out_word = 8'hCD;
		16'h967C: out_word = 8'hB4;
		16'h967D: out_word = 8'h30;
		16'h967E: out_word = 8'hCD;
		16'h967F: out_word = 8'h1E;
		16'h9680: out_word = 8'h31;
		16'h9681: out_word = 8'h30;
		16'h9682: out_word = 8'h26;
		16'h9683: out_word = 8'h1B;
		16'h9684: out_word = 8'h21;
		16'h9685: out_word = 8'h23;
		16'h9686: out_word = 8'h00;
		16'h9687: out_word = 8'h19;
		16'h9688: out_word = 8'hEB;
		16'h9689: out_word = 8'hC5;
		16'h968A: out_word = 8'h78;
		16'h968B: out_word = 8'hB9;
		16'h968C: out_word = 8'h28;
		16'h968D: out_word = 8'h0C;
		16'h968E: out_word = 8'hC5;
		16'h968F: out_word = 8'h01;
		16'h9690: out_word = 8'h23;
		16'h9691: out_word = 8'h00;
		16'h9692: out_word = 8'hED;
		16'h9693: out_word = 8'hB8;
		16'h9694: out_word = 8'hC1;
		16'h9695: out_word = 8'h78;
		16'h9696: out_word = 8'h0D;
		16'h9697: out_word = 8'hB9;
		16'h9698: out_word = 8'h38;
		16'h9699: out_word = 8'hF4;
		16'h969A: out_word = 8'hEB;
		16'h969B: out_word = 8'h13;
		16'h969C: out_word = 8'hC1;
		16'h969D: out_word = 8'hE1;
		16'h969E: out_word = 8'hCD;
		16'h969F: out_word = 8'h2C;
		16'h96A0: out_word = 8'h36;
		16'h96A1: out_word = 8'h01;
		16'h96A2: out_word = 8'h23;
		16'h96A3: out_word = 8'h00;
		16'h96A4: out_word = 8'hED;
		16'h96A5: out_word = 8'hB0;
		16'h96A6: out_word = 8'h37;
		16'h96A7: out_word = 8'hC1;
		16'h96A8: out_word = 8'hC9;
		16'h96A9: out_word = 8'hE1;
		16'h96AA: out_word = 8'hC1;
		16'h96AB: out_word = 8'hC9;
		16'h96AC: out_word = 8'hD5;
		16'h96AD: out_word = 8'h26;
		16'h96AE: out_word = 8'h00;
		16'h96AF: out_word = 8'h68;
		16'h96B0: out_word = 8'h19;
		16'h96B1: out_word = 8'h57;
		16'h96B2: out_word = 8'h78;
		16'h96B3: out_word = 8'h5E;
		16'h96B4: out_word = 8'h72;
		16'h96B5: out_word = 8'h53;
		16'h96B6: out_word = 8'h23;
		16'h96B7: out_word = 8'h3C;
		16'h96B8: out_word = 8'hFE;
		16'h96B9: out_word = 8'h20;
		16'h96BA: out_word = 8'h38;
		16'h96BB: out_word = 8'hF7;
		16'h96BC: out_word = 8'h7B;
		16'h96BD: out_word = 8'hFE;
		16'h96BE: out_word = 8'h00;
		16'h96BF: out_word = 8'hD1;
		16'h96C0: out_word = 8'hC9;
		16'h96C1: out_word = 8'hD5;
		16'h96C2: out_word = 8'h21;
		16'h96C3: out_word = 8'h20;
		16'h96C4: out_word = 8'h00;
		16'h96C5: out_word = 8'h19;
		16'h96C6: out_word = 8'hE5;
		16'h96C7: out_word = 8'h57;
		16'h96C8: out_word = 8'h3E;
		16'h96C9: out_word = 8'h1F;
		16'h96CA: out_word = 8'h18;
		16'h96CB: out_word = 8'h07;
		16'h96CC: out_word = 8'h5E;
		16'h96CD: out_word = 8'h72;
		16'h96CE: out_word = 8'h53;
		16'h96CF: out_word = 8'hB8;
		16'h96D0: out_word = 8'h28;
		16'h96D1: out_word = 8'h04;
		16'h96D2: out_word = 8'h3D;
		16'h96D3: out_word = 8'h2B;
		16'h96D4: out_word = 8'h18;
		16'h96D5: out_word = 8'hF6;
		16'h96D6: out_word = 8'h7B;
		16'h96D7: out_word = 8'hFE;
		16'h96D8: out_word = 8'h00;
		16'h96D9: out_word = 8'hE1;
		16'h96DA: out_word = 8'hD1;
		16'h96DB: out_word = 8'hC9;
		16'h96DC: out_word = 8'hB1;
		16'h96DD: out_word = 8'hC9;
		16'h96DE: out_word = 8'hBC;
		16'h96DF: out_word = 8'hBE;
		16'h96E0: out_word = 8'hC3;
		16'h96E1: out_word = 8'hAF;
		16'h96E2: out_word = 8'hB4;
		16'h96E3: out_word = 8'h93;
		16'h96E4: out_word = 8'h91;
		16'h96E5: out_word = 8'h92;
		16'h96E6: out_word = 8'h95;
		16'h96E7: out_word = 8'h98;
		16'h96E8: out_word = 8'h98;
		16'h96E9: out_word = 8'h98;
		16'h96EA: out_word = 8'h98;
		16'h96EB: out_word = 8'h98;
		16'h96EC: out_word = 8'h98;
		16'h96ED: out_word = 8'h98;
		16'h96EE: out_word = 8'h7F;
		16'h96EF: out_word = 8'h81;
		16'h96F0: out_word = 8'h2E;
		16'h96F1: out_word = 8'h6C;
		16'h96F2: out_word = 8'h6E;
		16'h96F3: out_word = 8'h70;
		16'h96F4: out_word = 8'h48;
		16'h96F5: out_word = 8'h94;
		16'h96F6: out_word = 8'h56;
		16'h96F7: out_word = 8'h3F;
		16'h96F8: out_word = 8'h41;
		16'h96F9: out_word = 8'h2B;
		16'h96FA: out_word = 8'h17;
		16'h96FB: out_word = 8'h1F;
		16'h96FC: out_word = 8'h37;
		16'h96FD: out_word = 8'h77;
		16'h96FE: out_word = 8'h44;
		16'h96FF: out_word = 8'h0F;
		16'h9700: out_word = 8'h59;
		16'h9701: out_word = 8'h2B;
		16'h9702: out_word = 8'h43;
		16'h9703: out_word = 8'h2D;
		16'h9704: out_word = 8'h51;
		16'h9705: out_word = 8'h3A;
		16'h9706: out_word = 8'h6D;
		16'h9707: out_word = 8'h42;
		16'h9708: out_word = 8'h0D;
		16'h9709: out_word = 8'h49;
		16'h970A: out_word = 8'h5C;
		16'h970B: out_word = 8'h44;
		16'h970C: out_word = 8'h15;
		16'h970D: out_word = 8'h5D;
		16'h970E: out_word = 8'h01;
		16'h970F: out_word = 8'h3D;
		16'h9710: out_word = 8'h02;
		16'h9711: out_word = 8'h06;
		16'h9712: out_word = 8'h00;
		16'h9713: out_word = 8'h67;
		16'h9714: out_word = 8'h1E;
		16'h9715: out_word = 8'h06;
		16'h9716: out_word = 8'hCB;
		16'h9717: out_word = 8'h0E;
		16'h9718: out_word = 8'h67;
		16'h9719: out_word = 8'h19;
		16'h971A: out_word = 8'h06;
		16'h971B: out_word = 8'h0C;
		16'h971C: out_word = 8'h53;
		16'h971D: out_word = 8'h1A;
		16'h971E: out_word = 8'h00;
		16'h971F: out_word = 8'hEE;
		16'h9720: out_word = 8'h1C;
		16'h9721: out_word = 8'h0C;
		16'h9722: out_word = 8'h6F;
		16'h9723: out_word = 8'h1A;
		16'h9724: out_word = 8'h04;
		16'h9725: out_word = 8'h3D;
		16'h9726: out_word = 8'h06;
		16'h9727: out_word = 8'hCC;
		16'h9728: out_word = 8'h06;
		16'h9729: out_word = 8'h0E;
		16'h972A: out_word = 8'h81;
		16'h972B: out_word = 8'h19;
		16'h972C: out_word = 8'h04;
		16'h972D: out_word = 8'h00;
		16'h972E: out_word = 8'hAB;
		16'h972F: out_word = 8'h1D;
		16'h9730: out_word = 8'h0E;
		16'h9731: out_word = 8'h78;
		16'h9732: out_word = 8'h21;
		16'h9733: out_word = 8'h0E;
		16'h9734: out_word = 8'h8C;
		16'h9735: out_word = 8'h21;
		16'h9736: out_word = 8'h0E;
		16'h9737: out_word = 8'hD5;
		16'h9738: out_word = 8'h21;
		16'h9739: out_word = 8'h0E;
		16'h973A: out_word = 8'h62;
		16'h973B: out_word = 8'h18;
		16'h973C: out_word = 8'h0C;
		16'h973D: out_word = 8'hAA;
		16'h973E: out_word = 8'h21;
		16'h973F: out_word = 8'h0D;
		16'h9740: out_word = 8'h02;
		16'h9741: out_word = 8'h1A;
		16'h9742: out_word = 8'h0E;
		16'h9743: out_word = 8'h75;
		16'h9744: out_word = 8'h1B;
		16'h9745: out_word = 8'h08;
		16'h9746: out_word = 8'h00;
		16'h9747: out_word = 8'h80;
		16'h9748: out_word = 8'h1E;
		16'h9749: out_word = 8'h03;
		16'h974A: out_word = 8'h4F;
		16'h974B: out_word = 8'h1E;
		16'h974C: out_word = 8'h00;
		16'h974D: out_word = 8'h5F;
		16'h974E: out_word = 8'h1E;
		16'h974F: out_word = 8'h0D;
		16'h9750: out_word = 8'h0D;
		16'h9751: out_word = 8'h1A;
		16'h9752: out_word = 8'h00;
		16'h9753: out_word = 8'h6B;
		16'h9754: out_word = 8'h0D;
		16'h9755: out_word = 8'h09;
		16'h9756: out_word = 8'h00;
		16'h9757: out_word = 8'hDC;
		16'h9758: out_word = 8'h22;
		16'h9759: out_word = 8'h06;
		16'h975A: out_word = 8'h00;
		16'h975B: out_word = 8'h3A;
		16'h975C: out_word = 8'h1F;
		16'h975D: out_word = 8'h0E;
		16'h975E: out_word = 8'hAB;
		16'h975F: out_word = 8'h19;
		16'h9760: out_word = 8'h0E;
		16'h9761: out_word = 8'hEB;
		16'h9762: out_word = 8'h19;
		16'h9763: out_word = 8'h03;
		16'h9764: out_word = 8'h42;
		16'h9765: out_word = 8'h1E;
		16'h9766: out_word = 8'h09;
		16'h9767: out_word = 8'h0E;
		16'h9768: out_word = 8'hBE;
		16'h9769: out_word = 8'h21;
		16'h976A: out_word = 8'h0C;
		16'h976B: out_word = 8'hA7;
		16'h976C: out_word = 8'h21;
		16'h976D: out_word = 8'h0E;
		16'h976E: out_word = 8'h74;
		16'h976F: out_word = 8'h21;
		16'h9770: out_word = 8'h0E;
		16'h9771: out_word = 8'h71;
		16'h9772: out_word = 8'h1B;
		16'h9773: out_word = 8'h0B;
		16'h9774: out_word = 8'h0B;
		16'h9775: out_word = 8'h0B;
		16'h9776: out_word = 8'h0B;
		16'h9777: out_word = 8'h08;
		16'h9778: out_word = 8'h00;
		16'h9779: out_word = 8'hF8;
		16'h977A: out_word = 8'h03;
		16'h977B: out_word = 8'h09;
		16'h977C: out_word = 8'h0E;
		16'h977D: out_word = 8'hAE;
		16'h977E: out_word = 8'h21;
		16'h977F: out_word = 8'h07;
		16'h9780: out_word = 8'h07;
		16'h9781: out_word = 8'h07;
		16'h9782: out_word = 8'h07;
		16'h9783: out_word = 8'h07;
		16'h9784: out_word = 8'h07;
		16'h9785: out_word = 8'h08;
		16'h9786: out_word = 8'h00;
		16'h9787: out_word = 8'h7A;
		16'h9788: out_word = 8'h1E;
		16'h9789: out_word = 8'h06;
		16'h978A: out_word = 8'h00;
		16'h978B: out_word = 8'h94;
		16'h978C: out_word = 8'h22;
		16'h978D: out_word = 8'h0E;
		16'h978E: out_word = 8'h8C;
		16'h978F: out_word = 8'h1A;
		16'h9790: out_word = 8'h06;
		16'h9791: out_word = 8'h2C;
		16'h9792: out_word = 8'h0A;
		16'h9793: out_word = 8'h00;
		16'h9794: out_word = 8'h36;
		16'h9795: out_word = 8'h17;
		16'h9796: out_word = 8'h06;
		16'h9797: out_word = 8'h00;
		16'h9798: out_word = 8'hE5;
		16'h9799: out_word = 8'h16;
		16'h979A: out_word = 8'h0E;
		16'h979B: out_word = 8'h41;
		16'h979C: out_word = 8'h06;
		16'h979D: out_word = 8'h0A;
		16'h979E: out_word = 8'h2C;
		16'h979F: out_word = 8'h0A;
		16'h97A0: out_word = 8'h0C;
		16'h97A1: out_word = 8'hF0;
		16'h97A2: out_word = 8'h1A;
		16'h97A3: out_word = 8'h0E;
		16'h97A4: out_word = 8'h0C;
		16'h97A5: out_word = 8'h1C;
		16'h97A6: out_word = 8'h0E;
		16'h97A7: out_word = 8'hE5;
		16'h97A8: out_word = 8'h1B;
		16'h97A9: out_word = 8'h0C;
		16'h97AA: out_word = 8'h2B;
		16'h97AB: out_word = 8'h1B;
		16'h97AC: out_word = 8'h0E;
		16'h97AD: out_word = 8'h17;
		16'h97AE: out_word = 8'h23;
		16'h97AF: out_word = 8'hFD;
		16'h97B0: out_word = 8'hCB;
		16'h97B1: out_word = 8'h01;
		16'h97B2: out_word = 8'hBE;
		16'h97B3: out_word = 8'hEF;
		16'h97B4: out_word = 8'hFB;
		16'h97B5: out_word = 8'h19;
		16'h97B6: out_word = 8'hAF;
		16'h97B7: out_word = 8'h32;
		16'h97B8: out_word = 8'h47;
		16'h97B9: out_word = 8'h5C;
		16'h97BA: out_word = 8'h3D;
		16'h97BB: out_word = 8'h32;
		16'h97BC: out_word = 8'h3A;
		16'h97BD: out_word = 8'h5C;
		16'h97BE: out_word = 8'h18;
		16'h97BF: out_word = 8'h01;
		16'h97C0: out_word = 8'hE7;
		16'h97C1: out_word = 8'hEF;
		16'h97C2: out_word = 8'hBF;
		16'h97C3: out_word = 8'h16;
		16'h97C4: out_word = 8'hFD;
		16'h97C5: out_word = 8'h34;
		16'h97C6: out_word = 8'h0D;
		16'h97C7: out_word = 8'hFA;
		16'h97C8: out_word = 8'h12;
		16'h97C9: out_word = 8'h19;
		16'h97CA: out_word = 8'hDF;
		16'h97CB: out_word = 8'h06;
		16'h97CC: out_word = 8'h00;
		16'h97CD: out_word = 8'hFE;
		16'h97CE: out_word = 8'h0D;
		16'h97CF: out_word = 8'hCA;
		16'h97D0: out_word = 8'h63;
		16'h97D1: out_word = 8'h18;
		16'h97D2: out_word = 8'hFE;
		16'h97D3: out_word = 8'h3A;
		16'h97D4: out_word = 8'h28;
		16'h97D5: out_word = 8'hEA;
		16'h97D6: out_word = 8'h21;
		16'h97D7: out_word = 8'h21;
		16'h97D8: out_word = 8'h18;
		16'h97D9: out_word = 8'hE5;
		16'h97DA: out_word = 8'h4F;
		16'h97DB: out_word = 8'hE7;
		16'h97DC: out_word = 8'h79;
		16'h97DD: out_word = 8'hD6;
		16'h97DE: out_word = 8'hCE;
		16'h97DF: out_word = 8'h30;
		16'h97E0: out_word = 8'h13;
		16'h97E1: out_word = 8'hC6;
		16'h97E2: out_word = 8'hCE;
		16'h97E3: out_word = 8'h21;
		16'h97E4: out_word = 8'hA9;
		16'h97E5: out_word = 8'h17;
		16'h97E6: out_word = 8'hFE;
		16'h97E7: out_word = 8'hA3;
		16'h97E8: out_word = 8'h28;
		16'h97E9: out_word = 8'h16;
		16'h97EA: out_word = 8'h21;
		16'h97EB: out_word = 8'hAC;
		16'h97EC: out_word = 8'h17;
		16'h97ED: out_word = 8'hFE;
		16'h97EE: out_word = 8'hA4;
		16'h97EF: out_word = 8'h28;
		16'h97F0: out_word = 8'h0F;
		16'h97F1: out_word = 8'hC3;
		16'h97F2: out_word = 8'h12;
		16'h97F3: out_word = 8'h19;
		16'h97F4: out_word = 8'h4F;
		16'h97F5: out_word = 8'h21;
		16'h97F6: out_word = 8'hDC;
		16'h97F7: out_word = 8'h16;
		16'h97F8: out_word = 8'h09;
		16'h97F9: out_word = 8'h4E;
		16'h97FA: out_word = 8'h09;
		16'h97FB: out_word = 8'h18;
		16'h97FC: out_word = 8'h03;
		16'h97FD: out_word = 8'h2A;
		16'h97FE: out_word = 8'h74;
		16'h97FF: out_word = 8'h5C;
		16'h9800: out_word = 8'h7E;
		16'h9801: out_word = 8'h23;
		16'h9802: out_word = 8'h22;
		16'h9803: out_word = 8'h74;
		16'h9804: out_word = 8'h5C;
		16'h9805: out_word = 8'h01;
		16'h9806: out_word = 8'hFD;
		16'h9807: out_word = 8'h17;
		16'h9808: out_word = 8'hC5;
		16'h9809: out_word = 8'h4F;
		16'h980A: out_word = 8'hFE;
		16'h980B: out_word = 8'h20;
		16'h980C: out_word = 8'h30;
		16'h980D: out_word = 8'h0C;
		16'h980E: out_word = 8'h21;
		16'h980F: out_word = 8'hB5;
		16'h9810: out_word = 8'h18;
		16'h9811: out_word = 8'h06;
		16'h9812: out_word = 8'h00;
		16'h9813: out_word = 8'h09;
		16'h9814: out_word = 8'h4E;
		16'h9815: out_word = 8'h09;
		16'h9816: out_word = 8'hE5;
		16'h9817: out_word = 8'hDF;
		16'h9818: out_word = 8'h05;
		16'h9819: out_word = 8'hC9;
		16'h981A: out_word = 8'hDF;
		16'h981B: out_word = 8'hB9;
		16'h981C: out_word = 8'hC2;
		16'h981D: out_word = 8'h12;
		16'h981E: out_word = 8'h19;
		16'h981F: out_word = 8'hE7;
		16'h9820: out_word = 8'hC9;
		16'h9821: out_word = 8'hCD;
		16'h9822: out_word = 8'hD6;
		16'h9823: out_word = 8'h05;
		16'h9824: out_word = 8'h38;
		16'h9825: out_word = 8'h04;
		16'h9826: out_word = 8'hCD;
		16'h9827: out_word = 8'hAC;
		16'h9828: out_word = 8'h05;
		16'h9829: out_word = 8'h14;
		16'h982A: out_word = 8'hFD;
		16'h982B: out_word = 8'hCB;
		16'h982C: out_word = 8'h0A;
		16'h982D: out_word = 8'h7E;
		16'h982E: out_word = 8'hC2;
		16'h982F: out_word = 8'hA8;
		16'h9830: out_word = 8'h18;
		16'h9831: out_word = 8'h2A;
		16'h9832: out_word = 8'h42;
		16'h9833: out_word = 8'h5C;
		16'h9834: out_word = 8'hCB;
		16'h9835: out_word = 8'h7C;
		16'h9836: out_word = 8'h28;
		16'h9837: out_word = 8'h14;
		16'h9838: out_word = 8'h21;
		16'h9839: out_word = 8'hFE;
		16'h983A: out_word = 8'hFF;
		16'h983B: out_word = 8'h22;
		16'h983C: out_word = 8'h45;
		16'h983D: out_word = 8'h5C;
		16'h983E: out_word = 8'h2A;
		16'h983F: out_word = 8'h61;
		16'h9840: out_word = 8'h5C;
		16'h9841: out_word = 8'h2B;
		16'h9842: out_word = 8'hED;
		16'h9843: out_word = 8'h5B;
		16'h9844: out_word = 8'h59;
		16'h9845: out_word = 8'h5C;
		16'h9846: out_word = 8'h1B;
		16'h9847: out_word = 8'h3A;
		16'h9848: out_word = 8'h44;
		16'h9849: out_word = 8'h5C;
		16'h984A: out_word = 8'h18;
		16'h984B: out_word = 8'h36;
		16'h984C: out_word = 8'hEF;
		16'h984D: out_word = 8'h6E;
		16'h984E: out_word = 8'h19;
		16'h984F: out_word = 8'h3A;
		16'h9850: out_word = 8'h44;
		16'h9851: out_word = 8'h5C;
		16'h9852: out_word = 8'h28;
		16'h9853: out_word = 8'h1C;
		16'h9854: out_word = 8'hA7;
		16'h9855: out_word = 8'h20;
		16'h9856: out_word = 8'h46;
		16'h9857: out_word = 8'h47;
		16'h9858: out_word = 8'h7E;
		16'h9859: out_word = 8'hE6;
		16'h985A: out_word = 8'hC0;
		16'h985B: out_word = 8'h78;
		16'h985C: out_word = 8'h28;
		16'h985D: out_word = 8'h12;
		16'h985E: out_word = 8'hCD;
		16'h985F: out_word = 8'hAC;
		16'h9860: out_word = 8'h05;
		16'h9861: out_word = 8'hFF;
		16'h9862: out_word = 8'hC1;
		16'h9863: out_word = 8'hFD;
		16'h9864: out_word = 8'hCB;
		16'h9865: out_word = 8'h01;
		16'h9866: out_word = 8'h7E;
		16'h9867: out_word = 8'hC8;
		16'h9868: out_word = 8'h2A;
		16'h9869: out_word = 8'h55;
		16'h986A: out_word = 8'h5C;
		16'h986B: out_word = 8'h3E;
		16'h986C: out_word = 8'hC0;
		16'h986D: out_word = 8'hA6;
		16'h986E: out_word = 8'hC0;
		16'h986F: out_word = 8'hAF;
		16'h9870: out_word = 8'hFE;
		16'h9871: out_word = 8'h01;
		16'h9872: out_word = 8'hCE;
		16'h9873: out_word = 8'h00;
		16'h9874: out_word = 8'h56;
		16'h9875: out_word = 8'h23;
		16'h9876: out_word = 8'h5E;
		16'h9877: out_word = 8'hED;
		16'h9878: out_word = 8'h53;
		16'h9879: out_word = 8'h45;
		16'h987A: out_word = 8'h5C;
		16'h987B: out_word = 8'h23;
		16'h987C: out_word = 8'h5E;
		16'h987D: out_word = 8'h23;
		16'h987E: out_word = 8'h56;
		16'h987F: out_word = 8'hEB;
		16'h9880: out_word = 8'h19;
		16'h9881: out_word = 8'h23;
		16'h9882: out_word = 8'h22;
		16'h9883: out_word = 8'h55;
		16'h9884: out_word = 8'h5C;
		16'h9885: out_word = 8'hEB;
		16'h9886: out_word = 8'h22;
		16'h9887: out_word = 8'h5D;
		16'h9888: out_word = 8'h5C;
		16'h9889: out_word = 8'h57;
		16'h988A: out_word = 8'h1E;
		16'h988B: out_word = 8'h00;
		16'h988C: out_word = 8'hFD;
		16'h988D: out_word = 8'h36;
		16'h988E: out_word = 8'h0A;
		16'h988F: out_word = 8'hFF;
		16'h9890: out_word = 8'h15;
		16'h9891: out_word = 8'hFD;
		16'h9892: out_word = 8'h72;
		16'h9893: out_word = 8'h0D;
		16'h9894: out_word = 8'hCA;
		16'h9895: out_word = 8'hC0;
		16'h9896: out_word = 8'h17;
		16'h9897: out_word = 8'h14;
		16'h9898: out_word = 8'hEF;
		16'h9899: out_word = 8'h8B;
		16'h989A: out_word = 8'h19;
		16'h989B: out_word = 8'h28;
		16'h989C: out_word = 8'h0B;
		16'h989D: out_word = 8'hCD;
		16'h989E: out_word = 8'hAC;
		16'h989F: out_word = 8'h05;
		16'h98A0: out_word = 8'h16;
		16'h98A1: out_word = 8'hFD;
		16'h98A2: out_word = 8'hCB;
		16'h98A3: out_word = 8'h01;
		16'h98A4: out_word = 8'h7E;
		16'h98A5: out_word = 8'hC0;
		16'h98A6: out_word = 8'hC1;
		16'h98A7: out_word = 8'hC1;
		16'h98A8: out_word = 8'hDF;
		16'h98A9: out_word = 8'hFE;
		16'h98AA: out_word = 8'h0D;
		16'h98AB: out_word = 8'h28;
		16'h98AC: out_word = 8'hB6;
		16'h98AD: out_word = 8'hFE;
		16'h98AE: out_word = 8'h3A;
		16'h98AF: out_word = 8'hCA;
		16'h98B0: out_word = 8'hC0;
		16'h98B1: out_word = 8'h17;
		16'h98B2: out_word = 8'hC3;
		16'h98B3: out_word = 8'h12;
		16'h98B4: out_word = 8'h19;
		16'h98B5: out_word = 8'h24;
		16'h98B6: out_word = 8'h43;
		16'h98B7: out_word = 8'h46;
		16'h98B8: out_word = 8'h1E;
		16'h98B9: out_word = 8'h4C;
		16'h98BA: out_word = 8'h20;
		16'h98BB: out_word = 8'h53;
		16'h98BC: out_word = 8'h5E;
		16'h98BD: out_word = 8'h4D;
		16'h98BE: out_word = 8'h86;
		16'h98BF: out_word = 8'h57;
		16'h98C0: out_word = 8'h88;
		16'h98C1: out_word = 8'h06;
		16'h98C2: out_word = 8'h02;
		16'h98C3: out_word = 8'h05;
		16'h98C4: out_word = 8'hEF;
		16'h98C5: out_word = 8'hDE;
		16'h98C6: out_word = 8'h1C;
		16'h98C7: out_word = 8'hBF;
		16'h98C8: out_word = 8'hC1;
		16'h98C9: out_word = 8'hCC;
		16'h98CA: out_word = 8'hA1;
		16'h98CB: out_word = 8'h18;
		16'h98CC: out_word = 8'hEB;
		16'h98CD: out_word = 8'h2A;
		16'h98CE: out_word = 8'h74;
		16'h98CF: out_word = 8'h5C;
		16'h98D0: out_word = 8'h4E;
		16'h98D1: out_word = 8'h23;
		16'h98D2: out_word = 8'h46;
		16'h98D3: out_word = 8'hEB;
		16'h98D4: out_word = 8'hC5;
		16'h98D5: out_word = 8'hC9;
		16'h98D6: out_word = 8'hEF;
		16'h98D7: out_word = 8'hDE;
		16'h98D8: out_word = 8'h1C;
		16'h98D9: out_word = 8'hBF;
		16'h98DA: out_word = 8'hC1;
		16'h98DB: out_word = 8'hCC;
		16'h98DC: out_word = 8'hA1;
		16'h98DD: out_word = 8'h18;
		16'h98DE: out_word = 8'hEB;
		16'h98DF: out_word = 8'h2A;
		16'h98E0: out_word = 8'h74;
		16'h98E1: out_word = 8'h5C;
		16'h98E2: out_word = 8'h4E;
		16'h98E3: out_word = 8'h23;
		16'h98E4: out_word = 8'h46;
		16'h98E5: out_word = 8'hEB;
		16'h98E6: out_word = 8'hE5;
		16'h98E7: out_word = 8'h21;
		16'h98E8: out_word = 8'hF8;
		16'h98E9: out_word = 8'h18;
		16'h98EA: out_word = 8'h22;
		16'h98EB: out_word = 8'h5A;
		16'h98EC: out_word = 8'h5B;
		16'h98ED: out_word = 8'h21;
		16'h98EE: out_word = 8'h14;
		16'h98EF: out_word = 8'h5B;
		16'h98F0: out_word = 8'hE3;
		16'h98F1: out_word = 8'hE5;
		16'h98F2: out_word = 8'h60;
		16'h98F3: out_word = 8'h69;
		16'h98F4: out_word = 8'hE3;
		16'h98F5: out_word = 8'hC3;
		16'h98F6: out_word = 8'h00;
		16'h98F7: out_word = 8'h5B;
		16'h98F8: out_word = 8'hC9;
		16'h98F9: out_word = 8'hEF;
		16'h98FA: out_word = 8'h1F;
		16'h98FB: out_word = 8'h1C;
		16'h98FC: out_word = 8'hC9;
		16'h98FD: out_word = 8'hC1;
		16'h98FE: out_word = 8'hEF;
		16'h98FF: out_word = 8'h56;
		16'h9900: out_word = 8'h1C;
		16'h9901: out_word = 8'hCD;
		16'h9902: out_word = 8'hA1;
		16'h9903: out_word = 8'h18;
		16'h9904: out_word = 8'hC9;
		16'h9905: out_word = 8'hEF;
		16'h9906: out_word = 8'h6C;
		16'h9907: out_word = 8'h1C;
		16'h9908: out_word = 8'hC9;
		16'h9909: out_word = 8'hE7;
		16'h990A: out_word = 8'hEF;
		16'h990B: out_word = 8'h7A;
		16'h990C: out_word = 8'h1C;
		16'h990D: out_word = 8'hC9;
		16'h990E: out_word = 8'hEF;
		16'h990F: out_word = 8'h82;
		16'h9910: out_word = 8'h1C;
		16'h9911: out_word = 8'hC9;
		16'h9912: out_word = 8'hCD;
		16'h9913: out_word = 8'hAC;
		16'h9914: out_word = 8'h05;
		16'h9915: out_word = 8'h0B;
		16'h9916: out_word = 8'hEF;
		16'h9917: out_word = 8'h8C;
		16'h9918: out_word = 8'h1C;
		16'h9919: out_word = 8'hC9;
		16'h991A: out_word = 8'hFD;
		16'h991B: out_word = 8'hCB;
		16'h991C: out_word = 8'h01;
		16'h991D: out_word = 8'h7E;
		16'h991E: out_word = 8'hFD;
		16'h991F: out_word = 8'hCB;
		16'h9920: out_word = 8'h02;
		16'h9921: out_word = 8'h86;
		16'h9922: out_word = 8'h28;
		16'h9923: out_word = 8'h03;
		16'h9924: out_word = 8'hEF;
		16'h9925: out_word = 8'h4D;
		16'h9926: out_word = 8'h0D;
		16'h9927: out_word = 8'hF1;
		16'h9928: out_word = 8'h3A;
		16'h9929: out_word = 8'h74;
		16'h992A: out_word = 8'h5C;
		16'h992B: out_word = 8'hD6;
		16'h992C: out_word = 8'hA7;
		16'h992D: out_word = 8'hEF;
		16'h992E: out_word = 8'hFC;
		16'h992F: out_word = 8'h21;
		16'h9930: out_word = 8'hCD;
		16'h9931: out_word = 8'hA1;
		16'h9932: out_word = 8'h18;
		16'h9933: out_word = 8'h2A;
		16'h9934: out_word = 8'h8F;
		16'h9935: out_word = 8'h5C;
		16'h9936: out_word = 8'h22;
		16'h9937: out_word = 8'h8D;
		16'h9938: out_word = 8'h5C;
		16'h9939: out_word = 8'h21;
		16'h993A: out_word = 8'h91;
		16'h993B: out_word = 8'h5C;
		16'h993C: out_word = 8'h7E;
		16'h993D: out_word = 8'h07;
		16'h993E: out_word = 8'hAE;
		16'h993F: out_word = 8'hE6;
		16'h9940: out_word = 8'hAA;
		16'h9941: out_word = 8'hAE;
		16'h9942: out_word = 8'h77;
		16'h9943: out_word = 8'hC9;
		16'h9944: out_word = 8'hEF;
		16'h9945: out_word = 8'hBE;
		16'h9946: out_word = 8'h1C;
		16'h9947: out_word = 8'hC9;
		16'h9948: out_word = 8'hF1;
		16'h9949: out_word = 8'h3A;
		16'h994A: out_word = 8'h66;
		16'h994B: out_word = 8'h5B;
		16'h994C: out_word = 8'hE6;
		16'h994D: out_word = 8'h0F;
		16'h994E: out_word = 8'h32;
		16'h994F: out_word = 8'h66;
		16'h9950: out_word = 8'h5B;
		16'h9951: out_word = 8'h3A;
		16'h9952: out_word = 8'h74;
		16'h9953: out_word = 8'h5C;
		16'h9954: out_word = 8'hD6;
		16'h9955: out_word = 8'h74;
		16'h9956: out_word = 8'h32;
		16'h9957: out_word = 8'h74;
		16'h9958: out_word = 8'h5C;
		16'h9959: out_word = 8'hCA;
		16'h995A: out_word = 8'hEB;
		16'h995B: out_word = 8'h11;
		16'h995C: out_word = 8'h3D;
		16'h995D: out_word = 8'hCA;
		16'h995E: out_word = 8'hF2;
		16'h995F: out_word = 8'h11;
		16'h9960: out_word = 8'h3D;
		16'h9961: out_word = 8'hCA;
		16'h9962: out_word = 8'hF9;
		16'h9963: out_word = 8'h11;
		16'h9964: out_word = 8'hC3;
		16'h9965: out_word = 8'h00;
		16'h9966: out_word = 8'h12;
		16'h9967: out_word = 8'hC1;
		16'h9968: out_word = 8'hFD;
		16'h9969: out_word = 8'hCB;
		16'h996A: out_word = 8'h01;
		16'h996B: out_word = 8'h7E;
		16'h996C: out_word = 8'h28;
		16'h996D: out_word = 8'h10;
		16'h996E: out_word = 8'h2A;
		16'h996F: out_word = 8'h65;
		16'h9970: out_word = 8'h5C;
		16'h9971: out_word = 8'h11;
		16'h9972: out_word = 8'hFB;
		16'h9973: out_word = 8'hFF;
		16'h9974: out_word = 8'h19;
		16'h9975: out_word = 8'h22;
		16'h9976: out_word = 8'h65;
		16'h9977: out_word = 8'h5C;
		16'h9978: out_word = 8'hEF;
		16'h9979: out_word = 8'hE9;
		16'h997A: out_word = 8'h34;
		16'h997B: out_word = 8'hDA;
		16'h997C: out_word = 8'h63;
		16'h997D: out_word = 8'h18;
		16'h997E: out_word = 8'hC3;
		16'h997F: out_word = 8'hC1;
		16'h9980: out_word = 8'h17;
		16'h9981: out_word = 8'hFE;
		16'h9982: out_word = 8'hCD;
		16'h9983: out_word = 8'h20;
		16'h9984: out_word = 8'h09;
		16'h9985: out_word = 8'hE7;
		16'h9986: out_word = 8'hCD;
		16'h9987: out_word = 8'h0E;
		16'h9988: out_word = 8'h19;
		16'h9989: out_word = 8'hCD;
		16'h998A: out_word = 8'hA1;
		16'h998B: out_word = 8'h18;
		16'h998C: out_word = 8'h18;
		16'h998D: out_word = 8'h18;
		16'h998E: out_word = 8'hCD;
		16'h998F: out_word = 8'hA1;
		16'h9990: out_word = 8'h18;
		16'h9991: out_word = 8'h2A;
		16'h9992: out_word = 8'h65;
		16'h9993: out_word = 8'h5C;
		16'h9994: out_word = 8'h36;
		16'h9995: out_word = 8'h00;
		16'h9996: out_word = 8'h23;
		16'h9997: out_word = 8'h36;
		16'h9998: out_word = 8'h00;
		16'h9999: out_word = 8'h23;
		16'h999A: out_word = 8'h36;
		16'h999B: out_word = 8'h01;
		16'h999C: out_word = 8'h23;
		16'h999D: out_word = 8'h36;
		16'h999E: out_word = 8'h00;
		16'h999F: out_word = 8'h23;
		16'h99A0: out_word = 8'h36;
		16'h99A1: out_word = 8'h00;
		16'h99A2: out_word = 8'h23;
		16'h99A3: out_word = 8'h22;
		16'h99A4: out_word = 8'h65;
		16'h99A5: out_word = 8'h5C;
		16'h99A6: out_word = 8'hEF;
		16'h99A7: out_word = 8'h16;
		16'h99A8: out_word = 8'h1D;
		16'h99A9: out_word = 8'hC9;
		16'h99AA: out_word = 8'hE7;
		16'h99AB: out_word = 8'hCD;
		16'h99AC: out_word = 8'hF9;
		16'h99AD: out_word = 8'h18;
		16'h99AE: out_word = 8'hFD;
		16'h99AF: out_word = 8'hCB;
		16'h99B0: out_word = 8'h01;
		16'h99B1: out_word = 8'h7E;
		16'h99B2: out_word = 8'h28;
		16'h99B3: out_word = 8'h2E;
		16'h99B4: out_word = 8'hDF;
		16'h99B5: out_word = 8'h22;
		16'h99B6: out_word = 8'h5F;
		16'h99B7: out_word = 8'h5C;
		16'h99B8: out_word = 8'h2A;
		16'h99B9: out_word = 8'h57;
		16'h99BA: out_word = 8'h5C;
		16'h99BB: out_word = 8'h7E;
		16'h99BC: out_word = 8'hFE;
		16'h99BD: out_word = 8'h2C;
		16'h99BE: out_word = 8'h28;
		16'h99BF: out_word = 8'h0B;
		16'h99C0: out_word = 8'h1E;
		16'h99C1: out_word = 8'hE4;
		16'h99C2: out_word = 8'hEF;
		16'h99C3: out_word = 8'h86;
		16'h99C4: out_word = 8'h1D;
		16'h99C5: out_word = 8'h30;
		16'h99C6: out_word = 8'h04;
		16'h99C7: out_word = 8'hCD;
		16'h99C8: out_word = 8'hAC;
		16'h99C9: out_word = 8'h05;
		16'h99CA: out_word = 8'h0D;
		16'h99CB: out_word = 8'h23;
		16'h99CC: out_word = 8'h22;
		16'h99CD: out_word = 8'h5D;
		16'h99CE: out_word = 8'h5C;
		16'h99CF: out_word = 8'h7E;
		16'h99D0: out_word = 8'hEF;
		16'h99D1: out_word = 8'h56;
		16'h99D2: out_word = 8'h1C;
		16'h99D3: out_word = 8'hDF;
		16'h99D4: out_word = 8'h22;
		16'h99D5: out_word = 8'h57;
		16'h99D6: out_word = 8'h5C;
		16'h99D7: out_word = 8'h2A;
		16'h99D8: out_word = 8'h5F;
		16'h99D9: out_word = 8'h5C;
		16'h99DA: out_word = 8'hFD;
		16'h99DB: out_word = 8'h36;
		16'h99DC: out_word = 8'h26;
		16'h99DD: out_word = 8'h00;
		16'h99DE: out_word = 8'h22;
		16'h99DF: out_word = 8'h5D;
		16'h99E0: out_word = 8'h5C;
		16'h99E1: out_word = 8'h7E;
		16'h99E2: out_word = 8'hDF;
		16'h99E3: out_word = 8'hFE;
		16'h99E4: out_word = 8'h2C;
		16'h99E5: out_word = 8'h28;
		16'h99E6: out_word = 8'hC3;
		16'h99E7: out_word = 8'hCD;
		16'h99E8: out_word = 8'hA1;
		16'h99E9: out_word = 8'h18;
		16'h99EA: out_word = 8'hC9;
		16'h99EB: out_word = 8'hFD;
		16'h99EC: out_word = 8'hCB;
		16'h99ED: out_word = 8'h01;
		16'h99EE: out_word = 8'h7E;
		16'h99EF: out_word = 8'h20;
		16'h99F0: out_word = 8'h0B;
		16'h99F1: out_word = 8'hEF;
		16'h99F2: out_word = 8'hFB;
		16'h99F3: out_word = 8'h24;
		16'h99F4: out_word = 8'hFE;
		16'h99F5: out_word = 8'h2C;
		16'h99F6: out_word = 8'hC4;
		16'h99F7: out_word = 8'hA1;
		16'h99F8: out_word = 8'h18;
		16'h99F9: out_word = 8'hE7;
		16'h99FA: out_word = 8'h18;
		16'h99FB: out_word = 8'hF5;
		16'h99FC: out_word = 8'h3E;
		16'h99FD: out_word = 8'hE4;
		16'h99FE: out_word = 8'hEF;
		16'h99FF: out_word = 8'h39;
		16'h9A00: out_word = 8'h1E;
		16'h9A01: out_word = 8'hC9;
		16'h9A02: out_word = 8'hEF;
		16'h9A03: out_word = 8'h67;
		16'h9A04: out_word = 8'h1E;
		16'h9A05: out_word = 8'h01;
		16'h9A06: out_word = 8'h00;
		16'h9A07: out_word = 8'h00;
		16'h9A08: out_word = 8'hEF;
		16'h9A09: out_word = 8'h45;
		16'h9A0A: out_word = 8'h1E;
		16'h9A0B: out_word = 8'h18;
		16'h9A0C: out_word = 8'h03;
		16'h9A0D: out_word = 8'hEF;
		16'h9A0E: out_word = 8'h99;
		16'h9A0F: out_word = 8'h1E;
		16'h9A10: out_word = 8'h78;
		16'h9A11: out_word = 8'hB1;
		16'h9A12: out_word = 8'h20;
		16'h9A13: out_word = 8'h04;
		16'h9A14: out_word = 8'hED;
		16'h9A15: out_word = 8'h4B;
		16'h9A16: out_word = 8'hB2;
		16'h9A17: out_word = 8'h5C;
		16'h9A18: out_word = 8'hC5;
		16'h9A19: out_word = 8'hED;
		16'h9A1A: out_word = 8'h5B;
		16'h9A1B: out_word = 8'h4B;
		16'h9A1C: out_word = 8'h5C;
		16'h9A1D: out_word = 8'h2A;
		16'h9A1E: out_word = 8'h59;
		16'h9A1F: out_word = 8'h5C;
		16'h9A20: out_word = 8'h2B;
		16'h9A21: out_word = 8'hEF;
		16'h9A22: out_word = 8'hE5;
		16'h9A23: out_word = 8'h19;
		16'h9A24: out_word = 8'hEF;
		16'h9A25: out_word = 8'h6B;
		16'h9A26: out_word = 8'h0D;
		16'h9A27: out_word = 8'h2A;
		16'h9A28: out_word = 8'h65;
		16'h9A29: out_word = 8'h5C;
		16'h9A2A: out_word = 8'h11;
		16'h9A2B: out_word = 8'h32;
		16'h9A2C: out_word = 8'h00;
		16'h9A2D: out_word = 8'h19;
		16'h9A2E: out_word = 8'hD1;
		16'h9A2F: out_word = 8'hED;
		16'h9A30: out_word = 8'h52;
		16'h9A31: out_word = 8'h30;
		16'h9A32: out_word = 8'h08;
		16'h9A33: out_word = 8'h2A;
		16'h9A34: out_word = 8'hB4;
		16'h9A35: out_word = 8'h5C;
		16'h9A36: out_word = 8'hA7;
		16'h9A37: out_word = 8'hED;
		16'h9A38: out_word = 8'h52;
		16'h9A39: out_word = 8'h30;
		16'h9A3A: out_word = 8'h04;
		16'h9A3B: out_word = 8'hCD;
		16'h9A3C: out_word = 8'hAC;
		16'h9A3D: out_word = 8'h05;
		16'h9A3E: out_word = 8'h15;
		16'h9A3F: out_word = 8'hED;
		16'h9A40: out_word = 8'h53;
		16'h9A41: out_word = 8'hB2;
		16'h9A42: out_word = 8'h5C;
		16'h9A43: out_word = 8'hD1;
		16'h9A44: out_word = 8'hE1;
		16'h9A45: out_word = 8'hC1;
		16'h9A46: out_word = 8'hED;
		16'h9A47: out_word = 8'h7B;
		16'h9A48: out_word = 8'hB2;
		16'h9A49: out_word = 8'h5C;
		16'h9A4A: out_word = 8'h33;
		16'h9A4B: out_word = 8'hC5;
		16'h9A4C: out_word = 8'hE5;
		16'h9A4D: out_word = 8'hED;
		16'h9A4E: out_word = 8'h73;
		16'h9A4F: out_word = 8'h3D;
		16'h9A50: out_word = 8'h5C;
		16'h9A51: out_word = 8'hD5;
		16'h9A52: out_word = 8'hC9;
		16'h9A53: out_word = 8'hD1;
		16'h9A54: out_word = 8'hFD;
		16'h9A55: out_word = 8'h66;
		16'h9A56: out_word = 8'h0D;
		16'h9A57: out_word = 8'h24;
		16'h9A58: out_word = 8'hE3;
		16'h9A59: out_word = 8'h33;
		16'h9A5A: out_word = 8'hED;
		16'h9A5B: out_word = 8'h4B;
		16'h9A5C: out_word = 8'h45;
		16'h9A5D: out_word = 8'h5C;
		16'h9A5E: out_word = 8'hC5;
		16'h9A5F: out_word = 8'hE5;
		16'h9A60: out_word = 8'hED;
		16'h9A61: out_word = 8'h73;
		16'h9A62: out_word = 8'h3D;
		16'h9A63: out_word = 8'h5C;
		16'h9A64: out_word = 8'hD5;
		16'h9A65: out_word = 8'hEF;
		16'h9A66: out_word = 8'h67;
		16'h9A67: out_word = 8'h1E;
		16'h9A68: out_word = 8'h01;
		16'h9A69: out_word = 8'h14;
		16'h9A6A: out_word = 8'h00;
		16'h9A6B: out_word = 8'hEF;
		16'h9A6C: out_word = 8'h05;
		16'h9A6D: out_word = 8'h1F;
		16'h9A6E: out_word = 8'hC9;
		16'h9A6F: out_word = 8'hC1;
		16'h9A70: out_word = 8'hE1;
		16'h9A71: out_word = 8'hD1;
		16'h9A72: out_word = 8'h7A;
		16'h9A73: out_word = 8'hFE;
		16'h9A74: out_word = 8'h3E;
		16'h9A75: out_word = 8'h28;
		16'h9A76: out_word = 8'h0F;
		16'h9A77: out_word = 8'h3B;
		16'h9A78: out_word = 8'hE3;
		16'h9A79: out_word = 8'hEB;
		16'h9A7A: out_word = 8'hED;
		16'h9A7B: out_word = 8'h73;
		16'h9A7C: out_word = 8'h3D;
		16'h9A7D: out_word = 8'h5C;
		16'h9A7E: out_word = 8'hC5;
		16'h9A7F: out_word = 8'h22;
		16'h9A80: out_word = 8'h42;
		16'h9A81: out_word = 8'h5C;
		16'h9A82: out_word = 8'hFD;
		16'h9A83: out_word = 8'h72;
		16'h9A84: out_word = 8'h0A;
		16'h9A85: out_word = 8'hC9;
		16'h9A86: out_word = 8'hD5;
		16'h9A87: out_word = 8'hE5;
		16'h9A88: out_word = 8'hCD;
		16'h9A89: out_word = 8'hAC;
		16'h9A8A: out_word = 8'h05;
		16'h9A8B: out_word = 8'h06;
		16'h9A8C: out_word = 8'hFD;
		16'h9A8D: out_word = 8'hCB;
		16'h9A8E: out_word = 8'h01;
		16'h9A8F: out_word = 8'h7E;
		16'h9A90: out_word = 8'h28;
		16'h9A91: out_word = 8'h05;
		16'h9A92: out_word = 8'h3E;
		16'h9A93: out_word = 8'hCE;
		16'h9A94: out_word = 8'hC3;
		16'h9A95: out_word = 8'hFE;
		16'h9A96: out_word = 8'h19;
		16'h9A97: out_word = 8'hFD;
		16'h9A98: out_word = 8'hCB;
		16'h9A99: out_word = 8'h01;
		16'h9A9A: out_word = 8'hF6;
		16'h9A9B: out_word = 8'hEF;
		16'h9A9C: out_word = 8'h8D;
		16'h9A9D: out_word = 8'h2C;
		16'h9A9E: out_word = 8'h30;
		16'h9A9F: out_word = 8'h16;
		16'h9AA0: out_word = 8'hE7;
		16'h9AA1: out_word = 8'hFE;
		16'h9AA2: out_word = 8'h24;
		16'h9AA3: out_word = 8'h20;
		16'h9AA4: out_word = 8'h05;
		16'h9AA5: out_word = 8'hFD;
		16'h9AA6: out_word = 8'hCB;
		16'h9AA7: out_word = 8'h01;
		16'h9AA8: out_word = 8'hB6;
		16'h9AA9: out_word = 8'hE7;
		16'h9AAA: out_word = 8'hFE;
		16'h9AAB: out_word = 8'h28;
		16'h9AAC: out_word = 8'h20;
		16'h9AAD: out_word = 8'h3C;
		16'h9AAE: out_word = 8'hE7;
		16'h9AAF: out_word = 8'hFE;
		16'h9AB0: out_word = 8'h29;
		16'h9AB1: out_word = 8'h28;
		16'h9AB2: out_word = 8'h20;
		16'h9AB3: out_word = 8'hEF;
		16'h9AB4: out_word = 8'h8D;
		16'h9AB5: out_word = 8'h2C;
		16'h9AB6: out_word = 8'hD2;
		16'h9AB7: out_word = 8'h12;
		16'h9AB8: out_word = 8'h19;
		16'h9AB9: out_word = 8'hEB;
		16'h9ABA: out_word = 8'hE7;
		16'h9ABB: out_word = 8'hFE;
		16'h9ABC: out_word = 8'h24;
		16'h9ABD: out_word = 8'h20;
		16'h9ABE: out_word = 8'h02;
		16'h9ABF: out_word = 8'hEB;
		16'h9AC0: out_word = 8'hE7;
		16'h9AC1: out_word = 8'hEB;
		16'h9AC2: out_word = 8'h01;
		16'h9AC3: out_word = 8'h06;
		16'h9AC4: out_word = 8'h00;
		16'h9AC5: out_word = 8'hEF;
		16'h9AC6: out_word = 8'h55;
		16'h9AC7: out_word = 8'h16;
		16'h9AC8: out_word = 8'h23;
		16'h9AC9: out_word = 8'h23;
		16'h9ACA: out_word = 8'h36;
		16'h9ACB: out_word = 8'h0E;
		16'h9ACC: out_word = 8'hFE;
		16'h9ACD: out_word = 8'h2C;
		16'h9ACE: out_word = 8'h20;
		16'h9ACF: out_word = 8'h03;
		16'h9AD0: out_word = 8'hE7;
		16'h9AD1: out_word = 8'h18;
		16'h9AD2: out_word = 8'hE0;
		16'h9AD3: out_word = 8'hFE;
		16'h9AD4: out_word = 8'h29;
		16'h9AD5: out_word = 8'h20;
		16'h9AD6: out_word = 8'h13;
		16'h9AD7: out_word = 8'hE7;
		16'h9AD8: out_word = 8'hFE;
		16'h9AD9: out_word = 8'h3D;
		16'h9ADA: out_word = 8'h20;
		16'h9ADB: out_word = 8'h0E;
		16'h9ADC: out_word = 8'hE7;
		16'h9ADD: out_word = 8'h3A;
		16'h9ADE: out_word = 8'h3B;
		16'h9ADF: out_word = 8'h5C;
		16'h9AE0: out_word = 8'hF5;
		16'h9AE1: out_word = 8'hEF;
		16'h9AE2: out_word = 8'hFB;
		16'h9AE3: out_word = 8'h24;
		16'h9AE4: out_word = 8'hF1;
		16'h9AE5: out_word = 8'hFD;
		16'h9AE6: out_word = 8'hAE;
		16'h9AE7: out_word = 8'h01;
		16'h9AE8: out_word = 8'hE6;
		16'h9AE9: out_word = 8'h40;
		16'h9AEA: out_word = 8'hC2;
		16'h9AEB: out_word = 8'h12;
		16'h9AEC: out_word = 8'h19;
		16'h9AED: out_word = 8'hCD;
		16'h9AEE: out_word = 8'hA1;
		16'h9AEF: out_word = 8'h18;
		16'h9AF0: out_word = 8'hC9;
		16'h9AF1: out_word = 8'h21;
		16'h9AF2: out_word = 8'h0E;
		16'h9AF3: out_word = 8'hEC;
		16'h9AF4: out_word = 8'h36;
		16'h9AF5: out_word = 8'hFF;
		16'h9AF6: out_word = 8'hCD;
		16'h9AF7: out_word = 8'h20;
		16'h9AF8: out_word = 8'h1F;
		16'h9AF9: out_word = 8'hEF;
		16'h9AFA: out_word = 8'hB0;
		16'h9AFB: out_word = 8'h16;
		16'h9AFC: out_word = 8'h2A;
		16'h9AFD: out_word = 8'h59;
		16'h9AFE: out_word = 8'h5C;
		16'h9AFF: out_word = 8'h01;
		16'h9B00: out_word = 8'h03;
		16'h9B01: out_word = 8'h00;
		16'h9B02: out_word = 8'hEF;
		16'h9B03: out_word = 8'h55;
		16'h9B04: out_word = 8'h16;
		16'h9B05: out_word = 8'h21;
		16'h9B06: out_word = 8'h6E;
		16'h9B07: out_word = 8'h1B;
		16'h9B08: out_word = 8'hED;
		16'h9B09: out_word = 8'h5B;
		16'h9B0A: out_word = 8'h59;
		16'h9B0B: out_word = 8'h5C;
		16'h9B0C: out_word = 8'h01;
		16'h9B0D: out_word = 8'h03;
		16'h9B0E: out_word = 8'h00;
		16'h9B0F: out_word = 8'hED;
		16'h9B10: out_word = 8'hB0;
		16'h9B11: out_word = 8'hCD;
		16'h9B12: out_word = 8'h6B;
		16'h9B13: out_word = 8'h02;
		16'h9B14: out_word = 8'hCD;
		16'h9B15: out_word = 8'h20;
		16'h9B16: out_word = 8'h1F;
		16'h9B17: out_word = 8'hEF;
		16'h9B18: out_word = 8'hB0;
		16'h9B19: out_word = 8'h16;
		16'h9B1A: out_word = 8'h2A;
		16'h9B1B: out_word = 8'h59;
		16'h9B1C: out_word = 8'h5C;
		16'h9B1D: out_word = 8'h01;
		16'h9B1E: out_word = 8'h01;
		16'h9B1F: out_word = 8'h00;
		16'h9B20: out_word = 8'hEF;
		16'h9B21: out_word = 8'h55;
		16'h9B22: out_word = 8'h16;
		16'h9B23: out_word = 8'h2A;
		16'h9B24: out_word = 8'h59;
		16'h9B25: out_word = 8'h5C;
		16'h9B26: out_word = 8'h36;
		16'h9B27: out_word = 8'hE1;
		16'h9B28: out_word = 8'hCD;
		16'h9B29: out_word = 8'h6B;
		16'h9B2A: out_word = 8'h02;
		16'h9B2B: out_word = 8'hCD;
		16'h9B2C: out_word = 8'h53;
		16'h9B2D: out_word = 8'h1B;
		16'h9B2E: out_word = 8'hED;
		16'h9B2F: out_word = 8'h7B;
		16'h9B30: out_word = 8'h3D;
		16'h9B31: out_word = 8'h5C;
		16'h9B32: out_word = 8'hE1;
		16'h9B33: out_word = 8'h21;
		16'h9B34: out_word = 8'h03;
		16'h9B35: out_word = 8'h13;
		16'h9B36: out_word = 8'hE5;
		16'h9B37: out_word = 8'h21;
		16'h9B38: out_word = 8'h13;
		16'h9B39: out_word = 8'h00;
		16'h9B3A: out_word = 8'hE5;
		16'h9B3B: out_word = 8'h21;
		16'h9B3C: out_word = 8'h08;
		16'h9B3D: out_word = 8'h00;
		16'h9B3E: out_word = 8'hE5;
		16'h9B3F: out_word = 8'h3E;
		16'h9B40: out_word = 8'h20;
		16'h9B41: out_word = 8'h32;
		16'h9B42: out_word = 8'h5C;
		16'h9B43: out_word = 8'h5B;
		16'h9B44: out_word = 8'hC3;
		16'h9B45: out_word = 8'h00;
		16'h9B46: out_word = 8'h5B;
		16'h9B47: out_word = 8'h21;
		16'h9B48: out_word = 8'h00;
		16'h9B49: out_word = 8'h00;
		16'h9B4A: out_word = 8'hE5;
		16'h9B4B: out_word = 8'h3E;
		16'h9B4C: out_word = 8'h20;
		16'h9B4D: out_word = 8'h32;
		16'h9B4E: out_word = 8'h5C;
		16'h9B4F: out_word = 8'h5B;
		16'h9B50: out_word = 8'hC3;
		16'h9B51: out_word = 8'h00;
		16'h9B52: out_word = 8'h5B;
		16'h9B53: out_word = 8'h2A;
		16'h9B54: out_word = 8'h4F;
		16'h9B55: out_word = 8'h5C;
		16'h9B56: out_word = 8'h11;
		16'h9B57: out_word = 8'h05;
		16'h9B58: out_word = 8'h00;
		16'h9B59: out_word = 8'h19;
		16'h9B5A: out_word = 8'h11;
		16'h9B5B: out_word = 8'h0A;
		16'h9B5C: out_word = 8'h00;
		16'h9B5D: out_word = 8'hEB;
		16'h9B5E: out_word = 8'h19;
		16'h9B5F: out_word = 8'hEB;
		16'h9B60: out_word = 8'h01;
		16'h9B61: out_word = 8'h04;
		16'h9B62: out_word = 8'h00;
		16'h9B63: out_word = 8'hED;
		16'h9B64: out_word = 8'hB0;
		16'h9B65: out_word = 8'hFD;
		16'h9B66: out_word = 8'hCB;
		16'h9B67: out_word = 8'h30;
		16'h9B68: out_word = 8'h9E;
		16'h9B69: out_word = 8'hFD;
		16'h9B6A: out_word = 8'hCB;
		16'h9B6B: out_word = 8'h01;
		16'h9B6C: out_word = 8'hA6;
		16'h9B6D: out_word = 8'hC9;
		16'h9B6E: out_word = 8'hEF;
		16'h9B6F: out_word = 8'h22;
		16'h9B70: out_word = 8'h22;
		16'h9B71: out_word = 8'h3E;
		16'h9B72: out_word = 8'h03;
		16'h9B73: out_word = 8'h18;
		16'h9B74: out_word = 8'h02;
		16'h9B75: out_word = 8'h3E;
		16'h9B76: out_word = 8'h02;
		16'h9B77: out_word = 8'hFD;
		16'h9B78: out_word = 8'h36;
		16'h9B79: out_word = 8'h02;
		16'h9B7A: out_word = 8'h00;
		16'h9B7B: out_word = 8'hEF;
		16'h9B7C: out_word = 8'h30;
		16'h9B7D: out_word = 8'h25;
		16'h9B7E: out_word = 8'h28;
		16'h9B7F: out_word = 8'h03;
		16'h9B80: out_word = 8'hEF;
		16'h9B81: out_word = 8'h01;
		16'h9B82: out_word = 8'h16;
		16'h9B83: out_word = 8'hEF;
		16'h9B84: out_word = 8'h18;
		16'h9B85: out_word = 8'h00;
		16'h9B86: out_word = 8'hEF;
		16'h9B87: out_word = 8'h70;
		16'h9B88: out_word = 8'h20;
		16'h9B89: out_word = 8'h38;
		16'h9B8A: out_word = 8'h18;
		16'h9B8B: out_word = 8'hEF;
		16'h9B8C: out_word = 8'h18;
		16'h9B8D: out_word = 8'h00;
		16'h9B8E: out_word = 8'hFE;
		16'h9B8F: out_word = 8'h3B;
		16'h9B90: out_word = 8'h28;
		16'h9B91: out_word = 8'h04;
		16'h9B92: out_word = 8'hFE;
		16'h9B93: out_word = 8'h2C;
		16'h9B94: out_word = 8'h20;
		16'h9B95: out_word = 8'h08;
		16'h9B96: out_word = 8'hEF;
		16'h9B97: out_word = 8'h20;
		16'h9B98: out_word = 8'h00;
		16'h9B99: out_word = 8'hCD;
		16'h9B9A: out_word = 8'h0E;
		16'h9B9B: out_word = 8'h19;
		16'h9B9C: out_word = 8'h18;
		16'h9B9D: out_word = 8'h08;
		16'h9B9E: out_word = 8'hEF;
		16'h9B9F: out_word = 8'hE6;
		16'h9BA0: out_word = 8'h1C;
		16'h9BA1: out_word = 8'h18;
		16'h9BA2: out_word = 8'h03;
		16'h9BA3: out_word = 8'hEF;
		16'h9BA4: out_word = 8'hDE;
		16'h9BA5: out_word = 8'h1C;
		16'h9BA6: out_word = 8'hCD;
		16'h9BA7: out_word = 8'hA1;
		16'h9BA8: out_word = 8'h18;
		16'h9BA9: out_word = 8'hEF;
		16'h9BAA: out_word = 8'h25;
		16'h9BAB: out_word = 8'h18;
		16'h9BAC: out_word = 8'hC9;
		16'h9BAD: out_word = 8'hED;
		16'h9BAE: out_word = 8'h73;
		16'h9BAF: out_word = 8'h81;
		16'h9BB0: out_word = 8'h5B;
		16'h9BB1: out_word = 8'h31;
		16'h9BB2: out_word = 8'hFF;
		16'h9BB3: out_word = 8'h5B;
		16'h9BB4: out_word = 8'hCD;
		16'h9BB5: out_word = 8'h97;
		16'h9BB6: out_word = 8'h1C;
		16'h9BB7: out_word = 8'hED;
		16'h9BB8: out_word = 8'h4B;
		16'h9BB9: out_word = 8'h72;
		16'h9BBA: out_word = 8'h5B;
		16'h9BBB: out_word = 8'h21;
		16'h9BBC: out_word = 8'hF7;
		16'h9BBD: out_word = 8'hFF;
		16'h9BBE: out_word = 8'hF6;
		16'h9BBF: out_word = 8'hFF;
		16'h9BC0: out_word = 8'hED;
		16'h9BC1: out_word = 8'h42;
		16'h9BC2: out_word = 8'hCD;
		16'h9BC3: out_word = 8'hF3;
		16'h9BC4: out_word = 8'h1C;
		16'h9BC5: out_word = 8'h01;
		16'h9BC6: out_word = 8'h09;
		16'h9BC7: out_word = 8'h00;
		16'h9BC8: out_word = 8'h21;
		16'h9BC9: out_word = 8'h71;
		16'h9BCA: out_word = 8'h5B;
		16'h9BCB: out_word = 8'hCD;
		16'h9BCC: out_word = 8'hAC;
		16'h9BCD: out_word = 8'h1D;
		16'h9BCE: out_word = 8'h2A;
		16'h9BCF: out_word = 8'h74;
		16'h9BD0: out_word = 8'h5B;
		16'h9BD1: out_word = 8'hED;
		16'h9BD2: out_word = 8'h4B;
		16'h9BD3: out_word = 8'h72;
		16'h9BD4: out_word = 8'h5B;
		16'h9BD5: out_word = 8'hCD;
		16'h9BD6: out_word = 8'hAC;
		16'h9BD7: out_word = 8'h1D;
		16'h9BD8: out_word = 8'hCD;
		16'h9BD9: out_word = 8'h56;
		16'h9BDA: out_word = 8'h1D;
		16'h9BDB: out_word = 8'h3E;
		16'h9BDC: out_word = 8'h05;
		16'h9BDD: out_word = 8'hCD;
		16'h9BDE: out_word = 8'h64;
		16'h9BDF: out_word = 8'h1C;
		16'h9BE0: out_word = 8'hED;
		16'h9BE1: out_word = 8'h7B;
		16'h9BE2: out_word = 8'h81;
		16'h9BE3: out_word = 8'h5B;
		16'h9BE4: out_word = 8'hC9;
		16'h9BE5: out_word = 8'hEF;
		16'h9BE6: out_word = 8'h18;
		16'h9BE7: out_word = 8'h00;
		16'h9BE8: out_word = 8'hFE;
		16'h9BE9: out_word = 8'h21;
		16'h9BEA: out_word = 8'hC2;
		16'h9BEB: out_word = 8'h12;
		16'h9BEC: out_word = 8'h19;
		16'h9BED: out_word = 8'hEF;
		16'h9BEE: out_word = 8'h20;
		16'h9BEF: out_word = 8'h00;
		16'h9BF0: out_word = 8'hCD;
		16'h9BF1: out_word = 8'hA1;
		16'h9BF2: out_word = 8'h18;
		16'h9BF3: out_word = 8'h3E;
		16'h9BF4: out_word = 8'h02;
		16'h9BF5: out_word = 8'hEF;
		16'h9BF6: out_word = 8'h01;
		16'h9BF7: out_word = 8'h16;
		16'h9BF8: out_word = 8'hED;
		16'h9BF9: out_word = 8'h73;
		16'h9BFA: out_word = 8'h81;
		16'h9BFB: out_word = 8'h5B;
		16'h9BFC: out_word = 8'h31;
		16'h9BFD: out_word = 8'hFF;
		16'h9BFE: out_word = 8'h5B;
		16'h9BFF: out_word = 8'hCD;
		16'h9C00: out_word = 8'hD2;
		16'h9C01: out_word = 8'h20;
		16'h9C02: out_word = 8'h3E;
		16'h9C03: out_word = 8'h05;
		16'h9C04: out_word = 8'hCD;
		16'h9C05: out_word = 8'h64;
		16'h9C06: out_word = 8'h1C;
		16'h9C07: out_word = 8'hED;
		16'h9C08: out_word = 8'h7B;
		16'h9C09: out_word = 8'h81;
		16'h9C0A: out_word = 8'h5B;
		16'h9C0B: out_word = 8'hC9;
		16'h9C0C: out_word = 8'hEF;
		16'h9C0D: out_word = 8'h18;
		16'h9C0E: out_word = 8'h00;
		16'h9C0F: out_word = 8'hFE;
		16'h9C10: out_word = 8'h21;
		16'h9C11: out_word = 8'hC2;
		16'h9C12: out_word = 8'h12;
		16'h9C13: out_word = 8'h19;
		16'h9C14: out_word = 8'hCD;
		16'h9C15: out_word = 8'h93;
		16'h9C16: out_word = 8'h13;
		16'h9C17: out_word = 8'hCD;
		16'h9C18: out_word = 8'hA1;
		16'h9C19: out_word = 8'h18;
		16'h9C1A: out_word = 8'hED;
		16'h9C1B: out_word = 8'h73;
		16'h9C1C: out_word = 8'h81;
		16'h9C1D: out_word = 8'h5B;
		16'h9C1E: out_word = 8'h31;
		16'h9C1F: out_word = 8'hFF;
		16'h9C20: out_word = 8'h5B;
		16'h9C21: out_word = 8'hCD;
		16'h9C22: out_word = 8'h5F;
		16'h9C23: out_word = 8'h1F;
		16'h9C24: out_word = 8'h3E;
		16'h9C25: out_word = 8'h05;
		16'h9C26: out_word = 8'hCD;
		16'h9C27: out_word = 8'h64;
		16'h9C28: out_word = 8'h1C;
		16'h9C29: out_word = 8'hED;
		16'h9C2A: out_word = 8'h7B;
		16'h9C2B: out_word = 8'h81;
		16'h9C2C: out_word = 8'h5B;
		16'h9C2D: out_word = 8'hC9;
		16'h9C2E: out_word = 8'hED;
		16'h9C2F: out_word = 8'h73;
		16'h9C30: out_word = 8'h81;
		16'h9C31: out_word = 8'h5B;
		16'h9C32: out_word = 8'h31;
		16'h9C33: out_word = 8'hFF;
		16'h9C34: out_word = 8'h5B;
		16'h9C35: out_word = 8'hCD;
		16'h9C36: out_word = 8'h35;
		16'h9C37: out_word = 8'h1D;
		16'h9C38: out_word = 8'h21;
		16'h9C39: out_word = 8'h71;
		16'h9C3A: out_word = 8'h5B;
		16'h9C3B: out_word = 8'h01;
		16'h9C3C: out_word = 8'h09;
		16'h9C3D: out_word = 8'h00;
		16'h9C3E: out_word = 8'hCD;
		16'h9C3F: out_word = 8'h37;
		16'h9C40: out_word = 8'h1E;
		16'h9C41: out_word = 8'h3E;
		16'h9C42: out_word = 8'h05;
		16'h9C43: out_word = 8'hCD;
		16'h9C44: out_word = 8'h64;
		16'h9C45: out_word = 8'h1C;
		16'h9C46: out_word = 8'hED;
		16'h9C47: out_word = 8'h7B;
		16'h9C48: out_word = 8'h81;
		16'h9C49: out_word = 8'h5B;
		16'h9C4A: out_word = 8'hC9;
		16'h9C4B: out_word = 8'hED;
		16'h9C4C: out_word = 8'h73;
		16'h9C4D: out_word = 8'h81;
		16'h9C4E: out_word = 8'h5B;
		16'h9C4F: out_word = 8'h31;
		16'h9C50: out_word = 8'hFF;
		16'h9C51: out_word = 8'h5B;
		16'h9C52: out_word = 8'h42;
		16'h9C53: out_word = 8'h4B;
		16'h9C54: out_word = 8'hCD;
		16'h9C55: out_word = 8'h37;
		16'h9C56: out_word = 8'h1E;
		16'h9C57: out_word = 8'hCD;
		16'h9C58: out_word = 8'h56;
		16'h9C59: out_word = 8'h1D;
		16'h9C5A: out_word = 8'h3E;
		16'h9C5B: out_word = 8'h05;
		16'h9C5C: out_word = 8'hCD;
		16'h9C5D: out_word = 8'h64;
		16'h9C5E: out_word = 8'h1C;
		16'h9C5F: out_word = 8'hED;
		16'h9C60: out_word = 8'h7B;
		16'h9C61: out_word = 8'h81;
		16'h9C62: out_word = 8'h5B;
		16'h9C63: out_word = 8'hC9;
		16'h9C64: out_word = 8'hE5;
		16'h9C65: out_word = 8'hC5;
		16'h9C66: out_word = 8'h21;
		16'h9C67: out_word = 8'h81;
		16'h9C68: out_word = 8'h1C;
		16'h9C69: out_word = 8'h06;
		16'h9C6A: out_word = 8'h00;
		16'h9C6B: out_word = 8'h4F;
		16'h9C6C: out_word = 8'h09;
		16'h9C6D: out_word = 8'h4E;
		16'h9C6E: out_word = 8'hF3;
		16'h9C6F: out_word = 8'h3A;
		16'h9C70: out_word = 8'h5C;
		16'h9C71: out_word = 8'h5B;
		16'h9C72: out_word = 8'hE6;
		16'h9C73: out_word = 8'hF8;
		16'h9C74: out_word = 8'hB1;
		16'h9C75: out_word = 8'h32;
		16'h9C76: out_word = 8'h5C;
		16'h9C77: out_word = 8'h5B;
		16'h9C78: out_word = 8'h01;
		16'h9C79: out_word = 8'hFD;
		16'h9C7A: out_word = 8'h7F;
		16'h9C7B: out_word = 8'hED;
		16'h9C7C: out_word = 8'h79;
		16'h9C7D: out_word = 8'hFB;
		16'h9C7E: out_word = 8'hC1;
		16'h9C7F: out_word = 8'hE1;
		16'h9C80: out_word = 8'hC9;
		16'h9C81: out_word = 8'h01;
		16'h9C82: out_word = 8'h03;
		16'h9C83: out_word = 8'h04;
		16'h9C84: out_word = 8'h06;
		16'h9C85: out_word = 8'h07;
		16'h9C86: out_word = 8'h00;
		16'h9C87: out_word = 8'h11;
		16'h9C88: out_word = 8'h67;
		16'h9C89: out_word = 8'h5B;
		16'h9C8A: out_word = 8'hDD;
		16'h9C8B: out_word = 8'hE5;
		16'h9C8C: out_word = 8'hE1;
		16'h9C8D: out_word = 8'h06;
		16'h9C8E: out_word = 8'h0A;
		16'h9C8F: out_word = 8'h1A;
		16'h9C90: out_word = 8'h13;
		16'h9C91: out_word = 8'hBE;
		16'h9C92: out_word = 8'h23;
		16'h9C93: out_word = 8'hC0;
		16'h9C94: out_word = 8'h10;
		16'h9C95: out_word = 8'hF9;
		16'h9C96: out_word = 8'hC9;
		16'h9C97: out_word = 8'hCD;
		16'h9C98: out_word = 8'h12;
		16'h9C99: out_word = 8'h1D;
		16'h9C9A: out_word = 8'h28;
		16'h9C9B: out_word = 8'h04;
		16'h9C9C: out_word = 8'hCD;
		16'h9C9D: out_word = 8'hAC;
		16'h9C9E: out_word = 8'h05;
		16'h9C9F: out_word = 8'h20;
		16'h9CA0: out_word = 8'hDD;
		16'h9CA1: out_word = 8'hE5;
		16'h9CA2: out_word = 8'h01;
		16'h9CA3: out_word = 8'hEC;
		16'h9CA4: out_word = 8'h3F;
		16'h9CA5: out_word = 8'hDD;
		16'h9CA6: out_word = 8'h09;
		16'h9CA7: out_word = 8'hDD;
		16'h9CA8: out_word = 8'hE1;
		16'h9CA9: out_word = 8'h30;
		16'h9CAA: out_word = 8'h63;
		16'h9CAB: out_word = 8'h21;
		16'h9CAC: out_word = 8'hEC;
		16'h9CAD: out_word = 8'hFF;
		16'h9CAE: out_word = 8'h3E;
		16'h9CAF: out_word = 8'hFF;
		16'h9CB0: out_word = 8'hCD;
		16'h9CB1: out_word = 8'hF3;
		16'h9CB2: out_word = 8'h1C;
		16'h9CB3: out_word = 8'h21;
		16'h9CB4: out_word = 8'h66;
		16'h9CB5: out_word = 8'h5B;
		16'h9CB6: out_word = 8'hCB;
		16'h9CB7: out_word = 8'hD6;
		16'h9CB8: out_word = 8'hDD;
		16'h9CB9: out_word = 8'hE5;
		16'h9CBA: out_word = 8'hD1;
		16'h9CBB: out_word = 8'h21;
		16'h9CBC: out_word = 8'h67;
		16'h9CBD: out_word = 8'h5B;
		16'h9CBE: out_word = 8'h01;
		16'h9CBF: out_word = 8'h0A;
		16'h9CC0: out_word = 8'h00;
		16'h9CC1: out_word = 8'hED;
		16'h9CC2: out_word = 8'hB0;
		16'h9CC3: out_word = 8'hDD;
		16'h9CC4: out_word = 8'hCB;
		16'h9CC5: out_word = 8'h13;
		16'h9CC6: out_word = 8'hC6;
		16'h9CC7: out_word = 8'hDD;
		16'h9CC8: out_word = 8'h7E;
		16'h9CC9: out_word = 8'h0A;
		16'h9CCA: out_word = 8'hDD;
		16'h9CCB: out_word = 8'h77;
		16'h9CCC: out_word = 8'h10;
		16'h9CCD: out_word = 8'hDD;
		16'h9CCE: out_word = 8'h7E;
		16'h9CCF: out_word = 8'h0B;
		16'h9CD0: out_word = 8'hDD;
		16'h9CD1: out_word = 8'h77;
		16'h9CD2: out_word = 8'h11;
		16'h9CD3: out_word = 8'hDD;
		16'h9CD4: out_word = 8'h7E;
		16'h9CD5: out_word = 8'h0C;
		16'h9CD6: out_word = 8'hDD;
		16'h9CD7: out_word = 8'h77;
		16'h9CD8: out_word = 8'h12;
		16'h9CD9: out_word = 8'hAF;
		16'h9CDA: out_word = 8'hDD;
		16'h9CDB: out_word = 8'h77;
		16'h9CDC: out_word = 8'h0D;
		16'h9CDD: out_word = 8'hDD;
		16'h9CDE: out_word = 8'h77;
		16'h9CDF: out_word = 8'h0E;
		16'h9CE0: out_word = 8'hDD;
		16'h9CE1: out_word = 8'h77;
		16'h9CE2: out_word = 8'h0F;
		16'h9CE3: out_word = 8'h3E;
		16'h9CE4: out_word = 8'h05;
		16'h9CE5: out_word = 8'hCD;
		16'h9CE6: out_word = 8'h64;
		16'h9CE7: out_word = 8'h1C;
		16'h9CE8: out_word = 8'hDD;
		16'h9CE9: out_word = 8'hE5;
		16'h9CEA: out_word = 8'hE1;
		16'h9CEB: out_word = 8'h01;
		16'h9CEC: out_word = 8'hEC;
		16'h9CED: out_word = 8'hFF;
		16'h9CEE: out_word = 8'h09;
		16'h9CEF: out_word = 8'h22;
		16'h9CF0: out_word = 8'h83;
		16'h9CF1: out_word = 8'h5B;
		16'h9CF2: out_word = 8'hC9;
		16'h9CF3: out_word = 8'hED;
		16'h9CF4: out_word = 8'h5B;
		16'h9CF5: out_word = 8'h85;
		16'h9CF6: out_word = 8'h5B;
		16'h9CF7: out_word = 8'h08;
		16'h9CF8: out_word = 8'h3A;
		16'h9CF9: out_word = 8'h87;
		16'h9CFA: out_word = 8'h5B;
		16'h9CFB: out_word = 8'h4F;
		16'h9CFC: out_word = 8'h08;
		16'h9CFD: out_word = 8'hCB;
		16'h9CFE: out_word = 8'h7F;
		16'h9CFF: out_word = 8'h20;
		16'h9D00: out_word = 8'h09;
		16'h9D01: out_word = 8'h19;
		16'h9D02: out_word = 8'h89;
		16'h9D03: out_word = 8'h22;
		16'h9D04: out_word = 8'h85;
		16'h9D05: out_word = 8'h5B;
		16'h9D06: out_word = 8'h32;
		16'h9D07: out_word = 8'h87;
		16'h9D08: out_word = 8'h5B;
		16'h9D09: out_word = 8'hC9;
		16'h9D0A: out_word = 8'h19;
		16'h9D0B: out_word = 8'h89;
		16'h9D0C: out_word = 8'h38;
		16'h9D0D: out_word = 8'hF5;
		16'h9D0E: out_word = 8'hCD;
		16'h9D0F: out_word = 8'hAC;
		16'h9D10: out_word = 8'h05;
		16'h9D11: out_word = 8'h03;
		16'h9D12: out_word = 8'h3E;
		16'h9D13: out_word = 8'h04;
		16'h9D14: out_word = 8'hCD;
		16'h9D15: out_word = 8'h64;
		16'h9D16: out_word = 8'h1C;
		16'h9D17: out_word = 8'hDD;
		16'h9D18: out_word = 8'h21;
		16'h9D19: out_word = 8'hEC;
		16'h9D1A: out_word = 8'hEB;
		16'h9D1B: out_word = 8'hED;
		16'h9D1C: out_word = 8'h5B;
		16'h9D1D: out_word = 8'h83;
		16'h9D1E: out_word = 8'h5B;
		16'h9D1F: out_word = 8'hB7;
		16'h9D20: out_word = 8'hDD;
		16'h9D21: out_word = 8'hE5;
		16'h9D22: out_word = 8'hE1;
		16'h9D23: out_word = 8'hED;
		16'h9D24: out_word = 8'h52;
		16'h9D25: out_word = 8'hC8;
		16'h9D26: out_word = 8'hCD;
		16'h9D27: out_word = 8'h87;
		16'h9D28: out_word = 8'h1C;
		16'h9D29: out_word = 8'h20;
		16'h9D2A: out_word = 8'h03;
		16'h9D2B: out_word = 8'hF6;
		16'h9D2C: out_word = 8'hFF;
		16'h9D2D: out_word = 8'hC9;
		16'h9D2E: out_word = 8'h01;
		16'h9D2F: out_word = 8'hEC;
		16'h9D30: out_word = 8'hFF;
		16'h9D31: out_word = 8'hDD;
		16'h9D32: out_word = 8'h09;
		16'h9D33: out_word = 8'h18;
		16'h9D34: out_word = 8'hE6;
		16'h9D35: out_word = 8'hCD;
		16'h9D36: out_word = 8'h12;
		16'h9D37: out_word = 8'h1D;
		16'h9D38: out_word = 8'h20;
		16'h9D39: out_word = 8'h04;
		16'h9D3A: out_word = 8'hCD;
		16'h9D3B: out_word = 8'hAC;
		16'h9D3C: out_word = 8'h05;
		16'h9D3D: out_word = 8'h23;
		16'h9D3E: out_word = 8'hDD;
		16'h9D3F: out_word = 8'h7E;
		16'h9D40: out_word = 8'h0A;
		16'h9D41: out_word = 8'hDD;
		16'h9D42: out_word = 8'h77;
		16'h9D43: out_word = 8'h10;
		16'h9D44: out_word = 8'hDD;
		16'h9D45: out_word = 8'h7E;
		16'h9D46: out_word = 8'h0B;
		16'h9D47: out_word = 8'hDD;
		16'h9D48: out_word = 8'h77;
		16'h9D49: out_word = 8'h11;
		16'h9D4A: out_word = 8'hDD;
		16'h9D4B: out_word = 8'h7E;
		16'h9D4C: out_word = 8'h0C;
		16'h9D4D: out_word = 8'hDD;
		16'h9D4E: out_word = 8'h77;
		16'h9D4F: out_word = 8'h12;
		16'h9D50: out_word = 8'h3E;
		16'h9D51: out_word = 8'h05;
		16'h9D52: out_word = 8'hCD;
		16'h9D53: out_word = 8'h64;
		16'h9D54: out_word = 8'h1C;
		16'h9D55: out_word = 8'hC9;
		16'h9D56: out_word = 8'h3E;
		16'h9D57: out_word = 8'h04;
		16'h9D58: out_word = 8'hCD;
		16'h9D59: out_word = 8'h64;
		16'h9D5A: out_word = 8'h1C;
		16'h9D5B: out_word = 8'hDD;
		16'h9D5C: out_word = 8'hCB;
		16'h9D5D: out_word = 8'h13;
		16'h9D5E: out_word = 8'h46;
		16'h9D5F: out_word = 8'hC8;
		16'h9D60: out_word = 8'hDD;
		16'h9D61: out_word = 8'hCB;
		16'h9D62: out_word = 8'h13;
		16'h9D63: out_word = 8'h86;
		16'h9D64: out_word = 8'h21;
		16'h9D65: out_word = 8'h66;
		16'h9D66: out_word = 8'h5B;
		16'h9D67: out_word = 8'hCB;
		16'h9D68: out_word = 8'h96;
		16'h9D69: out_word = 8'hDD;
		16'h9D6A: out_word = 8'h6E;
		16'h9D6B: out_word = 8'h10;
		16'h9D6C: out_word = 8'hDD;
		16'h9D6D: out_word = 8'h66;
		16'h9D6E: out_word = 8'h11;
		16'h9D6F: out_word = 8'hDD;
		16'h9D70: out_word = 8'h7E;
		16'h9D71: out_word = 8'h12;
		16'h9D72: out_word = 8'hDD;
		16'h9D73: out_word = 8'h5E;
		16'h9D74: out_word = 8'h0A;
		16'h9D75: out_word = 8'hDD;
		16'h9D76: out_word = 8'h56;
		16'h9D77: out_word = 8'h0B;
		16'h9D78: out_word = 8'hDD;
		16'h9D79: out_word = 8'h46;
		16'h9D7A: out_word = 8'h0C;
		16'h9D7B: out_word = 8'hB7;
		16'h9D7C: out_word = 8'hED;
		16'h9D7D: out_word = 8'h52;
		16'h9D7E: out_word = 8'h98;
		16'h9D7F: out_word = 8'hCB;
		16'h9D80: out_word = 8'h14;
		16'h9D81: out_word = 8'hCB;
		16'h9D82: out_word = 8'h14;
		16'h9D83: out_word = 8'hCB;
		16'h9D84: out_word = 8'h2F;
		16'h9D85: out_word = 8'hCB;
		16'h9D86: out_word = 8'h1C;
		16'h9D87: out_word = 8'hCB;
		16'h9D88: out_word = 8'h2F;
		16'h9D89: out_word = 8'hCB;
		16'h9D8A: out_word = 8'h1C;
		16'h9D8B: out_word = 8'hDD;
		16'h9D8C: out_word = 8'h75;
		16'h9D8D: out_word = 8'h0D;
		16'h9D8E: out_word = 8'hDD;
		16'h9D8F: out_word = 8'h74;
		16'h9D90: out_word = 8'h0E;
		16'h9D91: out_word = 8'hDD;
		16'h9D92: out_word = 8'h77;
		16'h9D93: out_word = 8'h0F;
		16'h9D94: out_word = 8'hDD;
		16'h9D95: out_word = 8'h6E;
		16'h9D96: out_word = 8'h10;
		16'h9D97: out_word = 8'hDD;
		16'h9D98: out_word = 8'h66;
		16'h9D99: out_word = 8'h11;
		16'h9D9A: out_word = 8'hDD;
		16'h9D9B: out_word = 8'h7E;
		16'h9D9C: out_word = 8'h12;
		16'h9D9D: out_word = 8'h01;
		16'h9D9E: out_word = 8'hEC;
		16'h9D9F: out_word = 8'hFF;
		16'h9DA0: out_word = 8'hDD;
		16'h9DA1: out_word = 8'h09;
		16'h9DA2: out_word = 8'hDD;
		16'h9DA3: out_word = 8'h75;
		16'h9DA4: out_word = 8'h0A;
		16'h9DA5: out_word = 8'hDD;
		16'h9DA6: out_word = 8'h74;
		16'h9DA7: out_word = 8'h0B;
		16'h9DA8: out_word = 8'hDD;
		16'h9DA9: out_word = 8'h77;
		16'h9DAA: out_word = 8'h0C;
		16'h9DAB: out_word = 8'hC9;
		16'h9DAC: out_word = 8'h78;
		16'h9DAD: out_word = 8'hB1;
		16'h9DAE: out_word = 8'hC8;
		16'h9DAF: out_word = 8'hE5;
		16'h9DB0: out_word = 8'h11;
		16'h9DB1: out_word = 8'h00;
		16'h9DB2: out_word = 8'hC0;
		16'h9DB3: out_word = 8'hEB;
		16'h9DB4: out_word = 8'hED;
		16'h9DB5: out_word = 8'h52;
		16'h9DB6: out_word = 8'h28;
		16'h9DB7: out_word = 8'h1D;
		16'h9DB8: out_word = 8'h38;
		16'h9DB9: out_word = 8'h1B;
		16'h9DBA: out_word = 8'hE5;
		16'h9DBB: out_word = 8'hED;
		16'h9DBC: out_word = 8'h42;
		16'h9DBD: out_word = 8'h30;
		16'h9DBE: out_word = 8'h0D;
		16'h9DBF: out_word = 8'h60;
		16'h9DC0: out_word = 8'h69;
		16'h9DC1: out_word = 8'hC1;
		16'h9DC2: out_word = 8'hB7;
		16'h9DC3: out_word = 8'hED;
		16'h9DC4: out_word = 8'h42;
		16'h9DC5: out_word = 8'hE3;
		16'h9DC6: out_word = 8'h11;
		16'h9DC7: out_word = 8'h00;
		16'h9DC8: out_word = 8'hC0;
		16'h9DC9: out_word = 8'hD5;
		16'h9DCA: out_word = 8'h18;
		16'h9DCB: out_word = 8'h28;
		16'h9DCC: out_word = 8'hE1;
		16'h9DCD: out_word = 8'hE1;
		16'h9DCE: out_word = 8'h11;
		16'h9DCF: out_word = 8'h00;
		16'h9DD0: out_word = 8'h00;
		16'h9DD1: out_word = 8'hD5;
		16'h9DD2: out_word = 8'hD5;
		16'h9DD3: out_word = 8'h18;
		16'h9DD4: out_word = 8'h1F;
		16'h9DD5: out_word = 8'h60;
		16'h9DD6: out_word = 8'h69;
		16'h9DD7: out_word = 8'h11;
		16'h9DD8: out_word = 8'h20;
		16'h9DD9: out_word = 8'h00;
		16'h9DDA: out_word = 8'hB7;
		16'h9DDB: out_word = 8'hED;
		16'h9DDC: out_word = 8'h52;
		16'h9DDD: out_word = 8'h38;
		16'h9DDE: out_word = 8'h05;
		16'h9DDF: out_word = 8'hE3;
		16'h9DE0: out_word = 8'h42;
		16'h9DE1: out_word = 8'h4B;
		16'h9DE2: out_word = 8'h18;
		16'h9DE3: out_word = 8'h05;
		16'h9DE4: out_word = 8'hE1;
		16'h9DE5: out_word = 8'h11;
		16'h9DE6: out_word = 8'h00;
		16'h9DE7: out_word = 8'h00;
		16'h9DE8: out_word = 8'hD5;
		16'h9DE9: out_word = 8'hC5;
		16'h9DEA: out_word = 8'h11;
		16'h9DEB: out_word = 8'h98;
		16'h9DEC: out_word = 8'h5B;
		16'h9DED: out_word = 8'hED;
		16'h9DEE: out_word = 8'hB0;
		16'h9DEF: out_word = 8'hC1;
		16'h9DF0: out_word = 8'hE5;
		16'h9DF1: out_word = 8'h21;
		16'h9DF2: out_word = 8'h98;
		16'h9DF3: out_word = 8'h5B;
		16'h9DF4: out_word = 8'h3E;
		16'h9DF5: out_word = 8'h04;
		16'h9DF6: out_word = 8'hCD;
		16'h9DF7: out_word = 8'h64;
		16'h9DF8: out_word = 8'h1C;
		16'h9DF9: out_word = 8'hDD;
		16'h9DFA: out_word = 8'h5E;
		16'h9DFB: out_word = 8'h10;
		16'h9DFC: out_word = 8'hDD;
		16'h9DFD: out_word = 8'h56;
		16'h9DFE: out_word = 8'h11;
		16'h9DFF: out_word = 8'hDD;
		16'h9E00: out_word = 8'h7E;
		16'h9E01: out_word = 8'h12;
		16'h9E02: out_word = 8'hCD;
		16'h9E03: out_word = 8'h64;
		16'h9E04: out_word = 8'h1C;
		16'h9E05: out_word = 8'hED;
		16'h9E06: out_word = 8'hA0;
		16'h9E07: out_word = 8'h7A;
		16'h9E08: out_word = 8'hB3;
		16'h9E09: out_word = 8'h28;
		16'h9E0A: out_word = 8'h19;
		16'h9E0B: out_word = 8'h78;
		16'h9E0C: out_word = 8'hB1;
		16'h9E0D: out_word = 8'hC2;
		16'h9E0E: out_word = 8'h05;
		16'h9E0F: out_word = 8'h1E;
		16'h9E10: out_word = 8'h3E;
		16'h9E11: out_word = 8'h04;
		16'h9E12: out_word = 8'hCD;
		16'h9E13: out_word = 8'h64;
		16'h9E14: out_word = 8'h1C;
		16'h9E15: out_word = 8'hDD;
		16'h9E16: out_word = 8'h73;
		16'h9E17: out_word = 8'h10;
		16'h9E18: out_word = 8'hDD;
		16'h9E19: out_word = 8'h72;
		16'h9E1A: out_word = 8'h11;
		16'h9E1B: out_word = 8'h3E;
		16'h9E1C: out_word = 8'h05;
		16'h9E1D: out_word = 8'hCD;
		16'h9E1E: out_word = 8'h64;
		16'h9E1F: out_word = 8'h1C;
		16'h9E20: out_word = 8'hE1;
		16'h9E21: out_word = 8'hC1;
		16'h9E22: out_word = 8'h18;
		16'h9E23: out_word = 8'h88;
		16'h9E24: out_word = 8'h3E;
		16'h9E25: out_word = 8'h04;
		16'h9E26: out_word = 8'hCD;
		16'h9E27: out_word = 8'h64;
		16'h9E28: out_word = 8'h1C;
		16'h9E29: out_word = 8'hDD;
		16'h9E2A: out_word = 8'h34;
		16'h9E2B: out_word = 8'h12;
		16'h9E2C: out_word = 8'hDD;
		16'h9E2D: out_word = 8'h7E;
		16'h9E2E: out_word = 8'h12;
		16'h9E2F: out_word = 8'h11;
		16'h9E30: out_word = 8'h00;
		16'h9E31: out_word = 8'hC0;
		16'h9E32: out_word = 8'hCD;
		16'h9E33: out_word = 8'h64;
		16'h9E34: out_word = 8'h1C;
		16'h9E35: out_word = 8'h18;
		16'h9E36: out_word = 8'hD4;
		16'h9E37: out_word = 8'h78;
		16'h9E38: out_word = 8'hB1;
		16'h9E39: out_word = 8'hC8;
		16'h9E3A: out_word = 8'hE5;
		16'h9E3B: out_word = 8'h11;
		16'h9E3C: out_word = 8'h00;
		16'h9E3D: out_word = 8'hC0;
		16'h9E3E: out_word = 8'hEB;
		16'h9E3F: out_word = 8'hED;
		16'h9E40: out_word = 8'h52;
		16'h9E41: out_word = 8'h28;
		16'h9E42: out_word = 8'h24;
		16'h9E43: out_word = 8'h38;
		16'h9E44: out_word = 8'h22;
		16'h9E45: out_word = 8'hE5;
		16'h9E46: out_word = 8'hED;
		16'h9E47: out_word = 8'h42;
		16'h9E48: out_word = 8'h30;
		16'h9E49: out_word = 8'h12;
		16'h9E4A: out_word = 8'h60;
		16'h9E4B: out_word = 8'h69;
		16'h9E4C: out_word = 8'hC1;
		16'h9E4D: out_word = 8'hB7;
		16'h9E4E: out_word = 8'hED;
		16'h9E4F: out_word = 8'h42;
		16'h9E50: out_word = 8'hE3;
		16'h9E51: out_word = 8'h11;
		16'h9E52: out_word = 8'h00;
		16'h9E53: out_word = 8'h00;
		16'h9E54: out_word = 8'hD5;
		16'h9E55: out_word = 8'h11;
		16'h9E56: out_word = 8'h00;
		16'h9E57: out_word = 8'hC0;
		16'h9E58: out_word = 8'hD5;
		16'h9E59: out_word = 8'hEB;
		16'h9E5A: out_word = 8'h18;
		16'h9E5B: out_word = 8'h24;
		16'h9E5C: out_word = 8'hE1;
		16'h9E5D: out_word = 8'hE1;
		16'h9E5E: out_word = 8'h11;
		16'h9E5F: out_word = 8'h00;
		16'h9E60: out_word = 8'h00;
		16'h9E61: out_word = 8'hD5;
		16'h9E62: out_word = 8'hD5;
		16'h9E63: out_word = 8'hD5;
		16'h9E64: out_word = 8'hEB;
		16'h9E65: out_word = 8'h18;
		16'h9E66: out_word = 8'h19;
		16'h9E67: out_word = 8'h60;
		16'h9E68: out_word = 8'h69;
		16'h9E69: out_word = 8'h11;
		16'h9E6A: out_word = 8'h20;
		16'h9E6B: out_word = 8'h00;
		16'h9E6C: out_word = 8'hB7;
		16'h9E6D: out_word = 8'hED;
		16'h9E6E: out_word = 8'h52;
		16'h9E6F: out_word = 8'h38;
		16'h9E70: out_word = 8'h05;
		16'h9E71: out_word = 8'hE3;
		16'h9E72: out_word = 8'h42;
		16'h9E73: out_word = 8'h4B;
		16'h9E74: out_word = 8'h18;
		16'h9E75: out_word = 8'h05;
		16'h9E76: out_word = 8'hE1;
		16'h9E77: out_word = 8'h11;
		16'h9E78: out_word = 8'h00;
		16'h9E79: out_word = 8'h00;
		16'h9E7A: out_word = 8'hD5;
		16'h9E7B: out_word = 8'hC5;
		16'h9E7C: out_word = 8'hE5;
		16'h9E7D: out_word = 8'h11;
		16'h9E7E: out_word = 8'h98;
		16'h9E7F: out_word = 8'h5B;
		16'h9E80: out_word = 8'h3E;
		16'h9E81: out_word = 8'h04;
		16'h9E82: out_word = 8'hCD;
		16'h9E83: out_word = 8'h64;
		16'h9E84: out_word = 8'h1C;
		16'h9E85: out_word = 8'hDD;
		16'h9E86: out_word = 8'h6E;
		16'h9E87: out_word = 8'h10;
		16'h9E88: out_word = 8'hDD;
		16'h9E89: out_word = 8'h66;
		16'h9E8A: out_word = 8'h11;
		16'h9E8B: out_word = 8'hDD;
		16'h9E8C: out_word = 8'h7E;
		16'h9E8D: out_word = 8'h12;
		16'h9E8E: out_word = 8'hCD;
		16'h9E8F: out_word = 8'h64;
		16'h9E90: out_word = 8'h1C;
		16'h9E91: out_word = 8'hED;
		16'h9E92: out_word = 8'hA0;
		16'h9E93: out_word = 8'h7C;
		16'h9E94: out_word = 8'hB5;
		16'h9E95: out_word = 8'h28;
		16'h9E96: out_word = 8'h25;
		16'h9E97: out_word = 8'h78;
		16'h9E98: out_word = 8'hB1;
		16'h9E99: out_word = 8'hC2;
		16'h9E9A: out_word = 8'h91;
		16'h9E9B: out_word = 8'h1E;
		16'h9E9C: out_word = 8'h3E;
		16'h9E9D: out_word = 8'h04;
		16'h9E9E: out_word = 8'hCD;
		16'h9E9F: out_word = 8'h64;
		16'h9EA0: out_word = 8'h1C;
		16'h9EA1: out_word = 8'hDD;
		16'h9EA2: out_word = 8'h75;
		16'h9EA3: out_word = 8'h10;
		16'h9EA4: out_word = 8'hDD;
		16'h9EA5: out_word = 8'h74;
		16'h9EA6: out_word = 8'h11;
		16'h9EA7: out_word = 8'h3E;
		16'h9EA8: out_word = 8'h05;
		16'h9EA9: out_word = 8'hCD;
		16'h9EAA: out_word = 8'h64;
		16'h9EAB: out_word = 8'h1C;
		16'h9EAC: out_word = 8'hD1;
		16'h9EAD: out_word = 8'hC1;
		16'h9EAE: out_word = 8'h21;
		16'h9EAF: out_word = 8'h98;
		16'h9EB0: out_word = 8'h5B;
		16'h9EB1: out_word = 8'h78;
		16'h9EB2: out_word = 8'hB1;
		16'h9EB3: out_word = 8'h28;
		16'h9EB4: out_word = 8'h02;
		16'h9EB5: out_word = 8'hED;
		16'h9EB6: out_word = 8'hB0;
		16'h9EB7: out_word = 8'hEB;
		16'h9EB8: out_word = 8'hC1;
		16'h9EB9: out_word = 8'hC3;
		16'h9EBA: out_word = 8'h37;
		16'h9EBB: out_word = 8'h1E;
		16'h9EBC: out_word = 8'h3E;
		16'h9EBD: out_word = 8'h04;
		16'h9EBE: out_word = 8'hCD;
		16'h9EBF: out_word = 8'h64;
		16'h9EC0: out_word = 8'h1C;
		16'h9EC1: out_word = 8'hDD;
		16'h9EC2: out_word = 8'h34;
		16'h9EC3: out_word = 8'h12;
		16'h9EC4: out_word = 8'hDD;
		16'h9EC5: out_word = 8'h7E;
		16'h9EC6: out_word = 8'h12;
		16'h9EC7: out_word = 8'h21;
		16'h9EC8: out_word = 8'h00;
		16'h9EC9: out_word = 8'hC0;
		16'h9ECA: out_word = 8'hCD;
		16'h9ECB: out_word = 8'h64;
		16'h9ECC: out_word = 8'h1C;
		16'h9ECD: out_word = 8'h18;
		16'h9ECE: out_word = 8'hC8;
		16'h9ECF: out_word = 8'hF5;
		16'h9ED0: out_word = 8'h3A;
		16'h9ED1: out_word = 8'h5C;
		16'h9ED2: out_word = 8'h5B;
		16'h9ED3: out_word = 8'hF5;
		16'h9ED4: out_word = 8'hE5;
		16'h9ED5: out_word = 8'hD5;
		16'h9ED6: out_word = 8'hC5;
		16'h9ED7: out_word = 8'hDD;
		16'h9ED8: out_word = 8'h21;
		16'h9ED9: out_word = 8'h6A;
		16'h9EDA: out_word = 8'h5B;
		16'h9EDB: out_word = 8'hDD;
		16'h9EDC: out_word = 8'h73;
		16'h9EDD: out_word = 8'h10;
		16'h9EDE: out_word = 8'hDD;
		16'h9EDF: out_word = 8'h72;
		16'h9EE0: out_word = 8'h11;
		16'h9EE1: out_word = 8'hDD;
		16'h9EE2: out_word = 8'h36;
		16'h9EE3: out_word = 8'h12;
		16'h9EE4: out_word = 8'h04;
		16'h9EE5: out_word = 8'hCD;
		16'h9EE6: out_word = 8'hAC;
		16'h9EE7: out_word = 8'h1D;
		16'h9EE8: out_word = 8'h3E;
		16'h9EE9: out_word = 8'h05;
		16'h9EEA: out_word = 8'hCD;
		16'h9EEB: out_word = 8'h64;
		16'h9EEC: out_word = 8'h1C;
		16'h9EED: out_word = 8'hC1;
		16'h9EEE: out_word = 8'hD1;
		16'h9EEF: out_word = 8'hE1;
		16'h9EF0: out_word = 8'h09;
		16'h9EF1: out_word = 8'hEB;
		16'h9EF2: out_word = 8'h09;
		16'h9EF3: out_word = 8'hEB;
		16'h9EF4: out_word = 8'hF1;
		16'h9EF5: out_word = 8'h01;
		16'h9EF6: out_word = 8'hFD;
		16'h9EF7: out_word = 8'h7F;
		16'h9EF8: out_word = 8'hF3;
		16'h9EF9: out_word = 8'hED;
		16'h9EFA: out_word = 8'h79;
		16'h9EFB: out_word = 8'h32;
		16'h9EFC: out_word = 8'h5C;
		16'h9EFD: out_word = 8'h5B;
		16'h9EFE: out_word = 8'hFB;
		16'h9EFF: out_word = 8'h01;
		16'h9F00: out_word = 8'h00;
		16'h9F01: out_word = 8'h00;
		16'h9F02: out_word = 8'hF1;
		16'h9F03: out_word = 8'hC9;
		16'h9F04: out_word = 8'hF5;
		16'h9F05: out_word = 8'h3A;
		16'h9F06: out_word = 8'h5C;
		16'h9F07: out_word = 8'h5B;
		16'h9F08: out_word = 8'hF5;
		16'h9F09: out_word = 8'hE5;
		16'h9F0A: out_word = 8'hD5;
		16'h9F0B: out_word = 8'hC5;
		16'h9F0C: out_word = 8'hDD;
		16'h9F0D: out_word = 8'h21;
		16'h9F0E: out_word = 8'h6A;
		16'h9F0F: out_word = 8'h5B;
		16'h9F10: out_word = 8'hDD;
		16'h9F11: out_word = 8'h75;
		16'h9F12: out_word = 8'h10;
		16'h9F13: out_word = 8'hDD;
		16'h9F14: out_word = 8'h74;
		16'h9F15: out_word = 8'h11;
		16'h9F16: out_word = 8'hDD;
		16'h9F17: out_word = 8'h36;
		16'h9F18: out_word = 8'h12;
		16'h9F19: out_word = 8'h04;
		16'h9F1A: out_word = 8'hEB;
		16'h9F1B: out_word = 8'hCD;
		16'h9F1C: out_word = 8'h37;
		16'h9F1D: out_word = 8'h1E;
		16'h9F1E: out_word = 8'h18;
		16'h9F1F: out_word = 8'hC8;
		16'h9F20: out_word = 8'h08;
		16'h9F21: out_word = 8'h3E;
		16'h9F22: out_word = 8'h00;
		16'h9F23: out_word = 8'hF3;
		16'h9F24: out_word = 8'hCD;
		16'h9F25: out_word = 8'h3A;
		16'h9F26: out_word = 8'h1F;
		16'h9F27: out_word = 8'hF1;
		16'h9F28: out_word = 8'h22;
		16'h9F29: out_word = 8'h58;
		16'h9F2A: out_word = 8'h5B;
		16'h9F2B: out_word = 8'h2A;
		16'h9F2C: out_word = 8'h81;
		16'h9F2D: out_word = 8'h5B;
		16'h9F2E: out_word = 8'hED;
		16'h9F2F: out_word = 8'h73;
		16'h9F30: out_word = 8'h81;
		16'h9F31: out_word = 8'h5B;
		16'h9F32: out_word = 8'hF9;
		16'h9F33: out_word = 8'hFB;
		16'h9F34: out_word = 8'h2A;
		16'h9F35: out_word = 8'h58;
		16'h9F36: out_word = 8'h5B;
		16'h9F37: out_word = 8'hF5;
		16'h9F38: out_word = 8'h08;
		16'h9F39: out_word = 8'hC9;
		16'h9F3A: out_word = 8'hC5;
		16'h9F3B: out_word = 8'h01;
		16'h9F3C: out_word = 8'hFD;
		16'h9F3D: out_word = 8'h7F;
		16'h9F3E: out_word = 8'hED;
		16'h9F3F: out_word = 8'h79;
		16'h9F40: out_word = 8'h32;
		16'h9F41: out_word = 8'h5C;
		16'h9F42: out_word = 8'h5B;
		16'h9F43: out_word = 8'hC1;
		16'h9F44: out_word = 8'hC9;
		16'h9F45: out_word = 8'h08;
		16'h9F46: out_word = 8'hF3;
		16'h9F47: out_word = 8'hF1;
		16'h9F48: out_word = 8'h22;
		16'h9F49: out_word = 8'h58;
		16'h9F4A: out_word = 8'h5B;
		16'h9F4B: out_word = 8'h2A;
		16'h9F4C: out_word = 8'h81;
		16'h9F4D: out_word = 8'h5B;
		16'h9F4E: out_word = 8'hED;
		16'h9F4F: out_word = 8'h73;
		16'h9F50: out_word = 8'h81;
		16'h9F51: out_word = 8'h5B;
		16'h9F52: out_word = 8'hF9;
		16'h9F53: out_word = 8'h2A;
		16'h9F54: out_word = 8'h58;
		16'h9F55: out_word = 8'h5B;
		16'h9F56: out_word = 8'hF5;
		16'h9F57: out_word = 8'h3E;
		16'h9F58: out_word = 8'h07;
		16'h9F59: out_word = 8'hCD;
		16'h9F5A: out_word = 8'h3A;
		16'h9F5B: out_word = 8'h1F;
		16'h9F5C: out_word = 8'hFB;
		16'h9F5D: out_word = 8'h08;
		16'h9F5E: out_word = 8'hC9;
		16'h9F5F: out_word = 8'hCD;
		16'h9F60: out_word = 8'h12;
		16'h9F61: out_word = 8'h1D;
		16'h9F62: out_word = 8'h20;
		16'h9F63: out_word = 8'h04;
		16'h9F64: out_word = 8'hCD;
		16'h9F65: out_word = 8'hAC;
		16'h9F66: out_word = 8'h05;
		16'h9F67: out_word = 8'h23;
		16'h9F68: out_word = 8'hDD;
		16'h9F69: out_word = 8'h6E;
		16'h9F6A: out_word = 8'h0D;
		16'h9F6B: out_word = 8'hDD;
		16'h9F6C: out_word = 8'h66;
		16'h9F6D: out_word = 8'h0E;
		16'h9F6E: out_word = 8'hDD;
		16'h9F6F: out_word = 8'h7E;
		16'h9F70: out_word = 8'h0F;
		16'h9F71: out_word = 8'hCD;
		16'h9F72: out_word = 8'hF3;
		16'h9F73: out_word = 8'h1C;
		16'h9F74: out_word = 8'hFD;
		16'h9F75: out_word = 8'hE5;
		16'h9F76: out_word = 8'hFD;
		16'h9F77: out_word = 8'h2A;
		16'h9F78: out_word = 8'h83;
		16'h9F79: out_word = 8'h5B;
		16'h9F7A: out_word = 8'h01;
		16'h9F7B: out_word = 8'hEC;
		16'h9F7C: out_word = 8'hFF;
		16'h9F7D: out_word = 8'hDD;
		16'h9F7E: out_word = 8'h09;
		16'h9F7F: out_word = 8'hFD;
		16'h9F80: out_word = 8'h6E;
		16'h9F81: out_word = 8'h0A;
		16'h9F82: out_word = 8'hFD;
		16'h9F83: out_word = 8'h66;
		16'h9F84: out_word = 8'h0B;
		16'h9F85: out_word = 8'hFD;
		16'h9F86: out_word = 8'h7E;
		16'h9F87: out_word = 8'h0C;
		16'h9F88: out_word = 8'hFD;
		16'h9F89: out_word = 8'hE1;
		16'h9F8A: out_word = 8'hDD;
		16'h9F8B: out_word = 8'h5E;
		16'h9F8C: out_word = 8'h0A;
		16'h9F8D: out_word = 8'hDD;
		16'h9F8E: out_word = 8'h56;
		16'h9F8F: out_word = 8'h0B;
		16'h9F90: out_word = 8'hDD;
		16'h9F91: out_word = 8'h46;
		16'h9F92: out_word = 8'h0C;
		16'h9F93: out_word = 8'hB7;
		16'h9F94: out_word = 8'hED;
		16'h9F95: out_word = 8'h52;
		16'h9F96: out_word = 8'h98;
		16'h9F97: out_word = 8'hCB;
		16'h9F98: out_word = 8'h14;
		16'h9F99: out_word = 8'hCB;
		16'h9F9A: out_word = 8'h14;
		16'h9F9B: out_word = 8'hCB;
		16'h9F9C: out_word = 8'h2F;
		16'h9F9D: out_word = 8'hCB;
		16'h9F9E: out_word = 8'h1C;
		16'h9F9F: out_word = 8'hCB;
		16'h9FA0: out_word = 8'h2F;
		16'h9FA1: out_word = 8'hCB;
		16'h9FA2: out_word = 8'h1C;
		16'h9FA3: out_word = 8'h01;
		16'h9FA4: out_word = 8'h14;
		16'h9FA5: out_word = 8'h00;
		16'h9FA6: out_word = 8'hDD;
		16'h9FA7: out_word = 8'h09;
		16'h9FA8: out_word = 8'hDD;
		16'h9FA9: out_word = 8'h75;
		16'h9FAA: out_word = 8'h10;
		16'h9FAB: out_word = 8'hDD;
		16'h9FAC: out_word = 8'h74;
		16'h9FAD: out_word = 8'h11;
		16'h9FAE: out_word = 8'hDD;
		16'h9FAF: out_word = 8'h77;
		16'h9FB0: out_word = 8'h12;
		16'h9FB1: out_word = 8'h01;
		16'h9FB2: out_word = 8'hEC;
		16'h9FB3: out_word = 8'hFF;
		16'h9FB4: out_word = 8'hDD;
		16'h9FB5: out_word = 8'h09;
		16'h9FB6: out_word = 8'hDD;
		16'h9FB7: out_word = 8'h6E;
		16'h9FB8: out_word = 8'h0A;
		16'h9FB9: out_word = 8'hDD;
		16'h9FBA: out_word = 8'h66;
		16'h9FBB: out_word = 8'h0B;
		16'h9FBC: out_word = 8'hDD;
		16'h9FBD: out_word = 8'h56;
		16'h9FBE: out_word = 8'h0C;
		16'h9FBF: out_word = 8'h01;
		16'h9FC0: out_word = 8'h14;
		16'h9FC1: out_word = 8'h00;
		16'h9FC2: out_word = 8'hDD;
		16'h9FC3: out_word = 8'h09;
		16'h9FC4: out_word = 8'h7A;
		16'h9FC5: out_word = 8'hCD;
		16'h9FC6: out_word = 8'h64;
		16'h9FC7: out_word = 8'h1C;
		16'h9FC8: out_word = 8'h3A;
		16'h9FC9: out_word = 8'h5C;
		16'h9FCA: out_word = 8'h5B;
		16'h9FCB: out_word = 8'h5F;
		16'h9FCC: out_word = 8'h01;
		16'h9FCD: out_word = 8'hFD;
		16'h9FCE: out_word = 8'h7F;
		16'h9FCF: out_word = 8'h3E;
		16'h9FD0: out_word = 8'h07;
		16'h9FD1: out_word = 8'hF3;
		16'h9FD2: out_word = 8'hED;
		16'h9FD3: out_word = 8'h79;
		16'h9FD4: out_word = 8'hD9;
		16'h9FD5: out_word = 8'hDD;
		16'h9FD6: out_word = 8'h6E;
		16'h9FD7: out_word = 8'h0A;
		16'h9FD8: out_word = 8'hDD;
		16'h9FD9: out_word = 8'h66;
		16'h9FDA: out_word = 8'h0B;
		16'h9FDB: out_word = 8'hDD;
		16'h9FDC: out_word = 8'h56;
		16'h9FDD: out_word = 8'h0C;
		16'h9FDE: out_word = 8'h7A;
		16'h9FDF: out_word = 8'hCD;
		16'h9FE0: out_word = 8'h64;
		16'h9FE1: out_word = 8'h1C;
		16'h9FE2: out_word = 8'h3A;
		16'h9FE3: out_word = 8'h5C;
		16'h9FE4: out_word = 8'h5B;
		16'h9FE5: out_word = 8'h5F;
		16'h9FE6: out_word = 8'h01;
		16'h9FE7: out_word = 8'hFD;
		16'h9FE8: out_word = 8'h7F;
		16'h9FE9: out_word = 8'hD9;
		16'h9FEA: out_word = 8'h3E;
		16'h9FEB: out_word = 8'h07;
		16'h9FEC: out_word = 8'hF3;
		16'h9FED: out_word = 8'hED;
		16'h9FEE: out_word = 8'h79;
		16'h9FEF: out_word = 8'hDD;
		16'h9FF0: out_word = 8'h7E;
		16'h9FF1: out_word = 8'h10;
		16'h9FF2: out_word = 8'hD6;
		16'h9FF3: out_word = 8'h01;
		16'h9FF4: out_word = 8'hDD;
		16'h9FF5: out_word = 8'h77;
		16'h9FF6: out_word = 8'h10;
		16'h9FF7: out_word = 8'h30;
		16'h9FF8: out_word = 8'h14;
		16'h9FF9: out_word = 8'hDD;
		16'h9FFA: out_word = 8'h7E;
		16'h9FFB: out_word = 8'h11;
		16'h9FFC: out_word = 8'hD6;
		16'h9FFD: out_word = 8'h01;
		16'h9FFE: out_word = 8'hDD;
		16'h9FFF: out_word = 8'h77;
		16'hA000: out_word = 8'h11;
		16'hA001: out_word = 8'h30;
		16'hA002: out_word = 8'h0A;
		16'hA003: out_word = 8'hDD;
		16'hA004: out_word = 8'h7E;
		16'hA005: out_word = 8'h12;
		16'hA006: out_word = 8'hD6;
		16'hA007: out_word = 8'h01;
		16'hA008: out_word = 8'hDD;
		16'hA009: out_word = 8'h77;
		16'hA00A: out_word = 8'h12;
		16'hA00B: out_word = 8'h38;
		16'hA00C: out_word = 8'h31;
		16'hA00D: out_word = 8'hED;
		16'hA00E: out_word = 8'h59;
		16'hA00F: out_word = 8'h7E;
		16'hA010: out_word = 8'h2C;
		16'hA011: out_word = 8'h20;
		16'hA012: out_word = 8'h11;
		16'hA013: out_word = 8'h24;
		16'hA014: out_word = 8'h20;
		16'hA015: out_word = 8'h0E;
		16'hA016: out_word = 8'h08;
		16'hA017: out_word = 8'h14;
		16'hA018: out_word = 8'h7A;
		16'hA019: out_word = 8'hCD;
		16'hA01A: out_word = 8'h64;
		16'hA01B: out_word = 8'h1C;
		16'hA01C: out_word = 8'h3A;
		16'hA01D: out_word = 8'h5C;
		16'hA01E: out_word = 8'h5B;
		16'hA01F: out_word = 8'h5F;
		16'hA020: out_word = 8'h21;
		16'hA021: out_word = 8'h00;
		16'hA022: out_word = 8'hC0;
		16'hA023: out_word = 8'h08;
		16'hA024: out_word = 8'hD9;
		16'hA025: out_word = 8'hF3;
		16'hA026: out_word = 8'hED;
		16'hA027: out_word = 8'h59;
		16'hA028: out_word = 8'h77;
		16'hA029: out_word = 8'h2C;
		16'hA02A: out_word = 8'h20;
		16'hA02B: out_word = 8'h0F;
		16'hA02C: out_word = 8'h24;
		16'hA02D: out_word = 8'h20;
		16'hA02E: out_word = 8'h0C;
		16'hA02F: out_word = 8'h14;
		16'hA030: out_word = 8'h7A;
		16'hA031: out_word = 8'hCD;
		16'hA032: out_word = 8'h64;
		16'hA033: out_word = 8'h1C;
		16'hA034: out_word = 8'h3A;
		16'hA035: out_word = 8'h5C;
		16'hA036: out_word = 8'h5B;
		16'hA037: out_word = 8'h5F;
		16'hA038: out_word = 8'h21;
		16'hA039: out_word = 8'h00;
		16'hA03A: out_word = 8'hC0;
		16'hA03B: out_word = 8'hD9;
		16'hA03C: out_word = 8'h18;
		16'hA03D: out_word = 8'hAC;
		16'hA03E: out_word = 8'h3E;
		16'hA03F: out_word = 8'h04;
		16'hA040: out_word = 8'hCD;
		16'hA041: out_word = 8'h64;
		16'hA042: out_word = 8'h1C;
		16'hA043: out_word = 8'h3E;
		16'hA044: out_word = 8'h00;
		16'hA045: out_word = 8'h21;
		16'hA046: out_word = 8'h14;
		16'hA047: out_word = 8'h00;
		16'hA048: out_word = 8'hCD;
		16'hA049: out_word = 8'hF3;
		16'hA04A: out_word = 8'h1C;
		16'hA04B: out_word = 8'hDD;
		16'hA04C: out_word = 8'h5E;
		16'hA04D: out_word = 8'h0D;
		16'hA04E: out_word = 8'hDD;
		16'hA04F: out_word = 8'h56;
		16'hA050: out_word = 8'h0E;
		16'hA051: out_word = 8'hDD;
		16'hA052: out_word = 8'h4E;
		16'hA053: out_word = 8'h0F;
		16'hA054: out_word = 8'h7A;
		16'hA055: out_word = 8'h07;
		16'hA056: out_word = 8'hCB;
		16'hA057: out_word = 8'h11;
		16'hA058: out_word = 8'h07;
		16'hA059: out_word = 8'hCB;
		16'hA05A: out_word = 8'h11;
		16'hA05B: out_word = 8'h7A;
		16'hA05C: out_word = 8'hE6;
		16'hA05D: out_word = 8'h3F;
		16'hA05E: out_word = 8'h57;
		16'hA05F: out_word = 8'hDD;
		16'hA060: out_word = 8'hE5;
		16'hA061: out_word = 8'hD5;
		16'hA062: out_word = 8'h11;
		16'hA063: out_word = 8'hEC;
		16'hA064: out_word = 8'hFF;
		16'hA065: out_word = 8'hDD;
		16'hA066: out_word = 8'h19;
		16'hA067: out_word = 8'hD1;
		16'hA068: out_word = 8'hDD;
		16'hA069: out_word = 8'h6E;
		16'hA06A: out_word = 8'h0A;
		16'hA06B: out_word = 8'hDD;
		16'hA06C: out_word = 8'h66;
		16'hA06D: out_word = 8'h0B;
		16'hA06E: out_word = 8'hDD;
		16'hA06F: out_word = 8'h7E;
		16'hA070: out_word = 8'h0C;
		16'hA071: out_word = 8'hB7;
		16'hA072: out_word = 8'hED;
		16'hA073: out_word = 8'h52;
		16'hA074: out_word = 8'h91;
		16'hA075: out_word = 8'hCB;
		16'hA076: out_word = 8'h74;
		16'hA077: out_word = 8'h20;
		16'hA078: out_word = 8'h03;
		16'hA079: out_word = 8'hCB;
		16'hA07A: out_word = 8'hF4;
		16'hA07B: out_word = 8'h3D;
		16'hA07C: out_word = 8'hDD;
		16'hA07D: out_word = 8'h75;
		16'hA07E: out_word = 8'h0A;
		16'hA07F: out_word = 8'hDD;
		16'hA080: out_word = 8'h74;
		16'hA081: out_word = 8'h0B;
		16'hA082: out_word = 8'hDD;
		16'hA083: out_word = 8'h77;
		16'hA084: out_word = 8'h0C;
		16'hA085: out_word = 8'hDD;
		16'hA086: out_word = 8'h6E;
		16'hA087: out_word = 8'h10;
		16'hA088: out_word = 8'hDD;
		16'hA089: out_word = 8'h66;
		16'hA08A: out_word = 8'h11;
		16'hA08B: out_word = 8'hDD;
		16'hA08C: out_word = 8'h7E;
		16'hA08D: out_word = 8'h12;
		16'hA08E: out_word = 8'hB7;
		16'hA08F: out_word = 8'hED;
		16'hA090: out_word = 8'h52;
		16'hA091: out_word = 8'h91;
		16'hA092: out_word = 8'hCB;
		16'hA093: out_word = 8'h74;
		16'hA094: out_word = 8'h20;
		16'hA095: out_word = 8'h03;
		16'hA096: out_word = 8'hCB;
		16'hA097: out_word = 8'hF4;
		16'hA098: out_word = 8'h3D;
		16'hA099: out_word = 8'hDD;
		16'hA09A: out_word = 8'h75;
		16'hA09B: out_word = 8'h10;
		16'hA09C: out_word = 8'hDD;
		16'hA09D: out_word = 8'h74;
		16'hA09E: out_word = 8'h11;
		16'hA09F: out_word = 8'hDD;
		16'hA0A0: out_word = 8'h77;
		16'hA0A1: out_word = 8'h12;
		16'hA0A2: out_word = 8'hDD;
		16'hA0A3: out_word = 8'hE5;
		16'hA0A4: out_word = 8'hE1;
		16'hA0A5: out_word = 8'hD5;
		16'hA0A6: out_word = 8'hED;
		16'hA0A7: out_word = 8'h5B;
		16'hA0A8: out_word = 8'h83;
		16'hA0A9: out_word = 8'h5B;
		16'hA0AA: out_word = 8'hB7;
		16'hA0AB: out_word = 8'hED;
		16'hA0AC: out_word = 8'h52;
		16'hA0AD: out_word = 8'hD1;
		16'hA0AE: out_word = 8'h20;
		16'hA0AF: out_word = 8'hB1;
		16'hA0B0: out_word = 8'hED;
		16'hA0B1: out_word = 8'h5B;
		16'hA0B2: out_word = 8'h83;
		16'hA0B3: out_word = 8'h5B;
		16'hA0B4: out_word = 8'hE1;
		16'hA0B5: out_word = 8'hE5;
		16'hA0B6: out_word = 8'hB7;
		16'hA0B7: out_word = 8'hED;
		16'hA0B8: out_word = 8'h52;
		16'hA0B9: out_word = 8'h44;
		16'hA0BA: out_word = 8'h4D;
		16'hA0BB: out_word = 8'hE1;
		16'hA0BC: out_word = 8'hE5;
		16'hA0BD: out_word = 8'h11;
		16'hA0BE: out_word = 8'h14;
		16'hA0BF: out_word = 8'h00;
		16'hA0C0: out_word = 8'h19;
		16'hA0C1: out_word = 8'hEB;
		16'hA0C2: out_word = 8'hE1;
		16'hA0C3: out_word = 8'h1B;
		16'hA0C4: out_word = 8'h2B;
		16'hA0C5: out_word = 8'hED;
		16'hA0C6: out_word = 8'hB8;
		16'hA0C7: out_word = 8'h2A;
		16'hA0C8: out_word = 8'h83;
		16'hA0C9: out_word = 8'h5B;
		16'hA0CA: out_word = 8'h11;
		16'hA0CB: out_word = 8'h14;
		16'hA0CC: out_word = 8'h00;
		16'hA0CD: out_word = 8'h19;
		16'hA0CE: out_word = 8'h22;
		16'hA0CF: out_word = 8'h83;
		16'hA0D0: out_word = 8'h5B;
		16'hA0D1: out_word = 8'hC9;
		16'hA0D2: out_word = 8'h3E;
		16'hA0D3: out_word = 8'h04;
		16'hA0D4: out_word = 8'hCD;
		16'hA0D5: out_word = 8'h64;
		16'hA0D6: out_word = 8'h1C;
		16'hA0D7: out_word = 8'h21;
		16'hA0D8: out_word = 8'h21;
		16'hA0D9: out_word = 8'h21;
		16'hA0DA: out_word = 8'h01;
		16'hA0DB: out_word = 8'h2B;
		16'hA0DC: out_word = 8'h21;
		16'hA0DD: out_word = 8'hDD;
		16'hA0DE: out_word = 8'h21;
		16'hA0DF: out_word = 8'hEC;
		16'hA0E0: out_word = 8'hEB;
		16'hA0E1: out_word = 8'hCD;
		16'hA0E2: out_word = 8'hD6;
		16'hA0E3: out_word = 8'h05;
		16'hA0E4: out_word = 8'hDD;
		16'hA0E5: out_word = 8'hE5;
		16'hA0E6: out_word = 8'hE3;
		16'hA0E7: out_word = 8'hED;
		16'hA0E8: out_word = 8'h5B;
		16'hA0E9: out_word = 8'h83;
		16'hA0EA: out_word = 8'h5B;
		16'hA0EB: out_word = 8'hB7;
		16'hA0EC: out_word = 8'hED;
		16'hA0ED: out_word = 8'h52;
		16'hA0EE: out_word = 8'hE1;
		16'hA0EF: out_word = 8'h28;
		16'hA0F0: out_word = 8'h20;
		16'hA0F1: out_word = 8'h54;
		16'hA0F2: out_word = 8'h5D;
		16'hA0F3: out_word = 8'hE5;
		16'hA0F4: out_word = 8'hC5;
		16'hA0F5: out_word = 8'hCD;
		16'hA0F6: out_word = 8'h8A;
		16'hA0F7: out_word = 8'h1C;
		16'hA0F8: out_word = 8'hC1;
		16'hA0F9: out_word = 8'hE1;
		16'hA0FA: out_word = 8'h30;
		16'hA0FB: out_word = 8'h0E;
		16'hA0FC: out_word = 8'h50;
		16'hA0FD: out_word = 8'h59;
		16'hA0FE: out_word = 8'hE5;
		16'hA0FF: out_word = 8'hC5;
		16'hA100: out_word = 8'hCD;
		16'hA101: out_word = 8'h8A;
		16'hA102: out_word = 8'h1C;
		16'hA103: out_word = 8'hC1;
		16'hA104: out_word = 8'hE1;
		16'hA105: out_word = 8'h38;
		16'hA106: out_word = 8'h03;
		16'hA107: out_word = 8'hDD;
		16'hA108: out_word = 8'hE5;
		16'hA109: out_word = 8'hC1;
		16'hA10A: out_word = 8'h11;
		16'hA10B: out_word = 8'hEC;
		16'hA10C: out_word = 8'hFF;
		16'hA10D: out_word = 8'hDD;
		16'hA10E: out_word = 8'h19;
		16'hA10F: out_word = 8'h18;
		16'hA110: out_word = 8'hD0;
		16'hA111: out_word = 8'hE5;
		16'hA112: out_word = 8'h21;
		16'hA113: out_word = 8'h2B;
		16'hA114: out_word = 8'h21;
		16'hA115: out_word = 8'hB7;
		16'hA116: out_word = 8'hED;
		16'hA117: out_word = 8'h42;
		16'hA118: out_word = 8'hE1;
		16'hA119: out_word = 8'hC8;
		16'hA11A: out_word = 8'h60;
		16'hA11B: out_word = 8'h69;
		16'hA11C: out_word = 8'hCD;
		16'hA11D: out_word = 8'h35;
		16'hA11E: out_word = 8'h21;
		16'hA11F: out_word = 8'h18;
		16'hA120: out_word = 8'hB9;
		16'hA121: out_word = 8'h00;
		16'hA122: out_word = 8'h00;
		16'hA123: out_word = 8'h00;
		16'hA124: out_word = 8'h00;
		16'hA125: out_word = 8'h00;
		16'hA126: out_word = 8'h00;
		16'hA127: out_word = 8'h00;
		16'hA128: out_word = 8'h00;
		16'hA129: out_word = 8'h00;
		16'hA12A: out_word = 8'h00;
		16'hA12B: out_word = 8'hFF;
		16'hA12C: out_word = 8'hFF;
		16'hA12D: out_word = 8'hFF;
		16'hA12E: out_word = 8'hFF;
		16'hA12F: out_word = 8'hFF;
		16'hA130: out_word = 8'hFF;
		16'hA131: out_word = 8'hFF;
		16'hA132: out_word = 8'hFF;
		16'hA133: out_word = 8'hFF;
		16'hA134: out_word = 8'hFF;
		16'hA135: out_word = 8'hE5;
		16'hA136: out_word = 8'hC5;
		16'hA137: out_word = 8'hE1;
		16'hA138: out_word = 8'h11;
		16'hA139: out_word = 8'h67;
		16'hA13A: out_word = 8'h5B;
		16'hA13B: out_word = 8'h01;
		16'hA13C: out_word = 8'h0A;
		16'hA13D: out_word = 8'h00;
		16'hA13E: out_word = 8'hED;
		16'hA13F: out_word = 8'hB0;
		16'hA140: out_word = 8'h3E;
		16'hA141: out_word = 8'h05;
		16'hA142: out_word = 8'hCD;
		16'hA143: out_word = 8'h64;
		16'hA144: out_word = 8'h1C;
		16'hA145: out_word = 8'h2A;
		16'hA146: out_word = 8'h81;
		16'hA147: out_word = 8'h5B;
		16'hA148: out_word = 8'hED;
		16'hA149: out_word = 8'h73;
		16'hA14A: out_word = 8'h81;
		16'hA14B: out_word = 8'h5B;
		16'hA14C: out_word = 8'hF9;
		16'hA14D: out_word = 8'h21;
		16'hA14E: out_word = 8'h67;
		16'hA14F: out_word = 8'h5B;
		16'hA150: out_word = 8'h06;
		16'hA151: out_word = 8'h0A;
		16'hA152: out_word = 8'h7E;
		16'hA153: out_word = 8'hE5;
		16'hA154: out_word = 8'hC5;
		16'hA155: out_word = 8'hEF;
		16'hA156: out_word = 8'h10;
		16'hA157: out_word = 8'h00;
		16'hA158: out_word = 8'hC1;
		16'hA159: out_word = 8'hE1;
		16'hA15A: out_word = 8'h23;
		16'hA15B: out_word = 8'h10;
		16'hA15C: out_word = 8'hF5;
		16'hA15D: out_word = 8'h3E;
		16'hA15E: out_word = 8'h0D;
		16'hA15F: out_word = 8'hEF;
		16'hA160: out_word = 8'h10;
		16'hA161: out_word = 8'h00;
		16'hA162: out_word = 8'hEF;
		16'hA163: out_word = 8'h4D;
		16'hA164: out_word = 8'h0D;
		16'hA165: out_word = 8'h2A;
		16'hA166: out_word = 8'h81;
		16'hA167: out_word = 8'h5B;
		16'hA168: out_word = 8'hED;
		16'hA169: out_word = 8'h73;
		16'hA16A: out_word = 8'h81;
		16'hA16B: out_word = 8'h5B;
		16'hA16C: out_word = 8'hF9;
		16'hA16D: out_word = 8'h3E;
		16'hA16E: out_word = 8'h04;
		16'hA16F: out_word = 8'hCD;
		16'hA170: out_word = 8'h64;
		16'hA171: out_word = 8'h1C;
		16'hA172: out_word = 8'hE1;
		16'hA173: out_word = 8'hC9;
		16'hA174: out_word = 8'h3E;
		16'hA175: out_word = 8'h03;
		16'hA176: out_word = 8'h18;
		16'hA177: out_word = 8'h02;
		16'hA178: out_word = 8'h3E;
		16'hA179: out_word = 8'h02;
		16'hA17A: out_word = 8'hEF;
		16'hA17B: out_word = 8'h30;
		16'hA17C: out_word = 8'h25;
		16'hA17D: out_word = 8'h28;
		16'hA17E: out_word = 8'h03;
		16'hA17F: out_word = 8'hEF;
		16'hA180: out_word = 8'h01;
		16'hA181: out_word = 8'h16;
		16'hA182: out_word = 8'hEF;
		16'hA183: out_word = 8'h4D;
		16'hA184: out_word = 8'h0D;
		16'hA185: out_word = 8'hEF;
		16'hA186: out_word = 8'hDF;
		16'hA187: out_word = 8'h1F;
		16'hA188: out_word = 8'hCD;
		16'hA189: out_word = 8'hA1;
		16'hA18A: out_word = 8'h18;
		16'hA18B: out_word = 8'hC9;
		16'hA18C: out_word = 8'hEF;
		16'hA18D: out_word = 8'h30;
		16'hA18E: out_word = 8'h25;
		16'hA18F: out_word = 8'h28;
		16'hA190: out_word = 8'h08;
		16'hA191: out_word = 8'h3E;
		16'hA192: out_word = 8'h01;
		16'hA193: out_word = 8'hEF;
		16'hA194: out_word = 8'h01;
		16'hA195: out_word = 8'h16;
		16'hA196: out_word = 8'hEF;
		16'hA197: out_word = 8'h6E;
		16'hA198: out_word = 8'h0D;
		16'hA199: out_word = 8'hFD;
		16'hA19A: out_word = 8'h36;
		16'hA19B: out_word = 8'h02;
		16'hA19C: out_word = 8'h01;
		16'hA19D: out_word = 8'hEF;
		16'hA19E: out_word = 8'hC1;
		16'hA19F: out_word = 8'h20;
		16'hA1A0: out_word = 8'hCD;
		16'hA1A1: out_word = 8'hA1;
		16'hA1A2: out_word = 8'h18;
		16'hA1A3: out_word = 8'hEF;
		16'hA1A4: out_word = 8'hA0;
		16'hA1A5: out_word = 8'h20;
		16'hA1A6: out_word = 8'hC9;
		16'hA1A7: out_word = 8'hC3;
		16'hA1A8: out_word = 8'hF0;
		16'hA1A9: out_word = 8'h08;
		16'hA1AA: out_word = 8'hF3;
		16'hA1AB: out_word = 8'hC3;
		16'hA1AC: out_word = 8'h9D;
		16'hA1AD: out_word = 8'h01;
		16'hA1AE: out_word = 8'hDF;
		16'hA1AF: out_word = 8'hFE;
		16'hA1B0: out_word = 8'h2C;
		16'hA1B1: out_word = 8'h20;
		16'hA1B2: out_word = 8'h38;
		16'hA1B3: out_word = 8'hE7;
		16'hA1B4: out_word = 8'hEF;
		16'hA1B5: out_word = 8'h82;
		16'hA1B6: out_word = 8'h1C;
		16'hA1B7: out_word = 8'hCD;
		16'hA1B8: out_word = 8'hA1;
		16'hA1B9: out_word = 8'h18;
		16'hA1BA: out_word = 8'hEF;
		16'hA1BB: out_word = 8'h2D;
		16'hA1BC: out_word = 8'h23;
		16'hA1BD: out_word = 8'hC9;
		16'hA1BE: out_word = 8'hDF;
		16'hA1BF: out_word = 8'hFE;
		16'hA1C0: out_word = 8'h2C;
		16'hA1C1: out_word = 8'h28;
		16'hA1C2: out_word = 8'h07;
		16'hA1C3: out_word = 8'hCD;
		16'hA1C4: out_word = 8'hA1;
		16'hA1C5: out_word = 8'h18;
		16'hA1C6: out_word = 8'hEF;
		16'hA1C7: out_word = 8'h77;
		16'hA1C8: out_word = 8'h24;
		16'hA1C9: out_word = 8'hC9;
		16'hA1CA: out_word = 8'hE7;
		16'hA1CB: out_word = 8'hEF;
		16'hA1CC: out_word = 8'h82;
		16'hA1CD: out_word = 8'h1C;
		16'hA1CE: out_word = 8'hCD;
		16'hA1CF: out_word = 8'hA1;
		16'hA1D0: out_word = 8'h18;
		16'hA1D1: out_word = 8'hEF;
		16'hA1D2: out_word = 8'h94;
		16'hA1D3: out_word = 8'h23;
		16'hA1D4: out_word = 8'hC9;
		16'hA1D5: out_word = 8'hEF;
		16'hA1D6: out_word = 8'hB2;
		16'hA1D7: out_word = 8'h28;
		16'hA1D8: out_word = 8'h20;
		16'hA1D9: out_word = 8'h11;
		16'hA1DA: out_word = 8'hEF;
		16'hA1DB: out_word = 8'h30;
		16'hA1DC: out_word = 8'h25;
		16'hA1DD: out_word = 8'h20;
		16'hA1DE: out_word = 8'h08;
		16'hA1DF: out_word = 8'hCB;
		16'hA1E0: out_word = 8'hB1;
		16'hA1E1: out_word = 8'hEF;
		16'hA1E2: out_word = 8'h96;
		16'hA1E3: out_word = 8'h29;
		16'hA1E4: out_word = 8'hCD;
		16'hA1E5: out_word = 8'hA1;
		16'hA1E6: out_word = 8'h18;
		16'hA1E7: out_word = 8'hEF;
		16'hA1E8: out_word = 8'h15;
		16'hA1E9: out_word = 8'h2C;
		16'hA1EA: out_word = 8'hC9;
		16'hA1EB: out_word = 8'hCD;
		16'hA1EC: out_word = 8'hAC;
		16'hA1ED: out_word = 8'h05;
		16'hA1EE: out_word = 8'h0B;
		16'hA1EF: out_word = 8'hFD;
		16'hA1F0: out_word = 8'hCB;
		16'hA1F1: out_word = 8'h30;
		16'hA1F2: out_word = 8'h46;
		16'hA1F3: out_word = 8'hC8;
		16'hA1F4: out_word = 8'hEF;
		16'hA1F5: out_word = 8'hAF;
		16'hA1F6: out_word = 8'h0D;
		16'hA1F7: out_word = 8'hC9;
		16'hA1F8: out_word = 8'h21;
		16'hA1F9: out_word = 8'hFE;
		16'hA1FA: out_word = 8'hFF;
		16'hA1FB: out_word = 8'h22;
		16'hA1FC: out_word = 8'h45;
		16'hA1FD: out_word = 8'h5C;
		16'hA1FE: out_word = 8'hFD;
		16'hA1FF: out_word = 8'hCB;
		16'hA200: out_word = 8'h01;
		16'hA201: out_word = 8'hBE;
		16'hA202: out_word = 8'hCD;
		16'hA203: out_word = 8'h8E;
		16'hA204: out_word = 8'h22;
		16'hA205: out_word = 8'hEF;
		16'hA206: out_word = 8'hFB;
		16'hA207: out_word = 8'h24;
		16'hA208: out_word = 8'hFD;
		16'hA209: out_word = 8'hCB;
		16'hA20A: out_word = 8'h01;
		16'hA20B: out_word = 8'h76;
		16'hA20C: out_word = 8'h28;
		16'hA20D: out_word = 8'h2C;
		16'hA20E: out_word = 8'hDF;
		16'hA20F: out_word = 8'hFE;
		16'hA210: out_word = 8'h0D;
		16'hA211: out_word = 8'h20;
		16'hA212: out_word = 8'h27;
		16'hA213: out_word = 8'hFD;
		16'hA214: out_word = 8'hCB;
		16'hA215: out_word = 8'h01;
		16'hA216: out_word = 8'hFE;
		16'hA217: out_word = 8'hCD;
		16'hA218: out_word = 8'h8E;
		16'hA219: out_word = 8'h22;
		16'hA21A: out_word = 8'h21;
		16'hA21B: out_word = 8'h21;
		16'hA21C: out_word = 8'h03;
		16'hA21D: out_word = 8'h22;
		16'hA21E: out_word = 8'h8B;
		16'hA21F: out_word = 8'h5B;
		16'hA220: out_word = 8'hEF;
		16'hA221: out_word = 8'hFB;
		16'hA222: out_word = 8'h24;
		16'hA223: out_word = 8'hFD;
		16'hA224: out_word = 8'hCB;
		16'hA225: out_word = 8'h01;
		16'hA226: out_word = 8'h76;
		16'hA227: out_word = 8'h28;
		16'hA228: out_word = 8'h11;
		16'hA229: out_word = 8'h11;
		16'hA22A: out_word = 8'h8D;
		16'hA22B: out_word = 8'h5B;
		16'hA22C: out_word = 8'h2A;
		16'hA22D: out_word = 8'h65;
		16'hA22E: out_word = 8'h5C;
		16'hA22F: out_word = 8'h01;
		16'hA230: out_word = 8'h05;
		16'hA231: out_word = 8'h00;
		16'hA232: out_word = 8'hB7;
		16'hA233: out_word = 8'hED;
		16'hA234: out_word = 8'h42;
		16'hA235: out_word = 8'hED;
		16'hA236: out_word = 8'hB0;
		16'hA237: out_word = 8'hC3;
		16'hA238: out_word = 8'h3E;
		16'hA239: out_word = 8'h22;
		16'hA23A: out_word = 8'hCD;
		16'hA23B: out_word = 8'hAC;
		16'hA23C: out_word = 8'h05;
		16'hA23D: out_word = 8'h19;
		16'hA23E: out_word = 8'h3E;
		16'hA23F: out_word = 8'h0D;
		16'hA240: out_word = 8'hCD;
		16'hA241: out_word = 8'h6F;
		16'hA242: out_word = 8'h22;
		16'hA243: out_word = 8'h01;
		16'hA244: out_word = 8'h01;
		16'hA245: out_word = 8'h00;
		16'hA246: out_word = 8'hEF;
		16'hA247: out_word = 8'h30;
		16'hA248: out_word = 8'h00;
		16'hA249: out_word = 8'h22;
		16'hA24A: out_word = 8'h5B;
		16'hA24B: out_word = 8'h5C;
		16'hA24C: out_word = 8'hE5;
		16'hA24D: out_word = 8'h2A;
		16'hA24E: out_word = 8'h51;
		16'hA24F: out_word = 8'h5C;
		16'hA250: out_word = 8'hE5;
		16'hA251: out_word = 8'h3E;
		16'hA252: out_word = 8'hFF;
		16'hA253: out_word = 8'hEF;
		16'hA254: out_word = 8'h01;
		16'hA255: out_word = 8'h16;
		16'hA256: out_word = 8'hEF;
		16'hA257: out_word = 8'hE3;
		16'hA258: out_word = 8'h2D;
		16'hA259: out_word = 8'hE1;
		16'hA25A: out_word = 8'hEF;
		16'hA25B: out_word = 8'h15;
		16'hA25C: out_word = 8'h16;
		16'hA25D: out_word = 8'hD1;
		16'hA25E: out_word = 8'h2A;
		16'hA25F: out_word = 8'h5B;
		16'hA260: out_word = 8'h5C;
		16'hA261: out_word = 8'hA7;
		16'hA262: out_word = 8'hED;
		16'hA263: out_word = 8'h52;
		16'hA264: out_word = 8'h1A;
		16'hA265: out_word = 8'hCD;
		16'hA266: out_word = 8'h6F;
		16'hA267: out_word = 8'h22;
		16'hA268: out_word = 8'h13;
		16'hA269: out_word = 8'h2B;
		16'hA26A: out_word = 8'h7C;
		16'hA26B: out_word = 8'hB5;
		16'hA26C: out_word = 8'h20;
		16'hA26D: out_word = 8'hF6;
		16'hA26E: out_word = 8'hC9;
		16'hA26F: out_word = 8'hE5;
		16'hA270: out_word = 8'hD5;
		16'hA271: out_word = 8'hCD;
		16'hA272: out_word = 8'h45;
		16'hA273: out_word = 8'h1F;
		16'hA274: out_word = 8'h21;
		16'hA275: out_word = 8'h0D;
		16'hA276: out_word = 8'hEC;
		16'hA277: out_word = 8'hCB;
		16'hA278: out_word = 8'h9E;
		16'hA279: out_word = 8'hF5;
		16'hA27A: out_word = 8'h3E;
		16'hA27B: out_word = 8'h02;
		16'hA27C: out_word = 8'hEF;
		16'hA27D: out_word = 8'h01;
		16'hA27E: out_word = 8'h16;
		16'hA27F: out_word = 8'hF1;
		16'hA280: out_word = 8'hCD;
		16'hA281: out_word = 8'h69;
		16'hA282: out_word = 8'h26;
		16'hA283: out_word = 8'h21;
		16'hA284: out_word = 8'h0D;
		16'hA285: out_word = 8'hEC;
		16'hA286: out_word = 8'hCB;
		16'hA287: out_word = 8'h9E;
		16'hA288: out_word = 8'hCD;
		16'hA289: out_word = 8'h20;
		16'hA28A: out_word = 8'h1F;
		16'hA28B: out_word = 8'hD1;
		16'hA28C: out_word = 8'hE1;
		16'hA28D: out_word = 8'hC9;
		16'hA28E: out_word = 8'h2A;
		16'hA28F: out_word = 8'h59;
		16'hA290: out_word = 8'h5C;
		16'hA291: out_word = 8'h2B;
		16'hA292: out_word = 8'h22;
		16'hA293: out_word = 8'h5D;
		16'hA294: out_word = 8'h5C;
		16'hA295: out_word = 8'hE7;
		16'hA296: out_word = 8'hC9;
		16'hA297: out_word = 8'hCD;
		16'hA298: out_word = 8'h8E;
		16'hA299: out_word = 8'h22;
		16'hA29A: out_word = 8'hFE;
		16'hA29B: out_word = 8'hF1;
		16'hA29C: out_word = 8'hC0;
		16'hA29D: out_word = 8'h2A;
		16'hA29E: out_word = 8'h5D;
		16'hA29F: out_word = 8'h5C;
		16'hA2A0: out_word = 8'h7E;
		16'hA2A1: out_word = 8'h23;
		16'hA2A2: out_word = 8'hFE;
		16'hA2A3: out_word = 8'h0D;
		16'hA2A4: out_word = 8'hC8;
		16'hA2A5: out_word = 8'hFE;
		16'hA2A6: out_word = 8'h3A;
		16'hA2A7: out_word = 8'h20;
		16'hA2A8: out_word = 8'hF7;
		16'hA2A9: out_word = 8'hB7;
		16'hA2AA: out_word = 8'hC9;
		16'hA2AB: out_word = 8'h47;
		16'hA2AC: out_word = 8'h21;
		16'hA2AD: out_word = 8'hBD;
		16'hA2AE: out_word = 8'h22;
		16'hA2AF: out_word = 8'h7E;
		16'hA2B0: out_word = 8'h23;
		16'hA2B1: out_word = 8'hB7;
		16'hA2B2: out_word = 8'h28;
		16'hA2B3: out_word = 8'h05;
		16'hA2B4: out_word = 8'hB8;
		16'hA2B5: out_word = 8'h20;
		16'hA2B6: out_word = 8'hF8;
		16'hA2B7: out_word = 8'h78;
		16'hA2B8: out_word = 8'hC9;
		16'hA2B9: out_word = 8'hF6;
		16'hA2BA: out_word = 8'hFF;
		16'hA2BB: out_word = 8'h78;
		16'hA2BC: out_word = 8'hC9;
		16'hA2BD: out_word = 8'h2B;
		16'hA2BE: out_word = 8'h2D;
		16'hA2BF: out_word = 8'h2A;
		16'hA2C0: out_word = 8'h2F;
		16'hA2C1: out_word = 8'h5E;
		16'hA2C2: out_word = 8'h3D;
		16'hA2C3: out_word = 8'h3E;
		16'hA2C4: out_word = 8'h3C;
		16'hA2C5: out_word = 8'hC7;
		16'hA2C6: out_word = 8'hC8;
		16'hA2C7: out_word = 8'hC9;
		16'hA2C8: out_word = 8'hC5;
		16'hA2C9: out_word = 8'hC6;
		16'hA2CA: out_word = 8'h00;
		16'hA2CB: out_word = 8'hFE;
		16'hA2CC: out_word = 8'hA5;
		16'hA2CD: out_word = 8'h38;
		16'hA2CE: out_word = 8'h0E;
		16'hA2CF: out_word = 8'hFE;
		16'hA2D0: out_word = 8'hC4;
		16'hA2D1: out_word = 8'h30;
		16'hA2D2: out_word = 8'h0A;
		16'hA2D3: out_word = 8'hFE;
		16'hA2D4: out_word = 8'hAC;
		16'hA2D5: out_word = 8'h28;
		16'hA2D6: out_word = 8'h06;
		16'hA2D7: out_word = 8'hFE;
		16'hA2D8: out_word = 8'hAD;
		16'hA2D9: out_word = 8'h28;
		16'hA2DA: out_word = 8'h02;
		16'hA2DB: out_word = 8'hBF;
		16'hA2DC: out_word = 8'hC9;
		16'hA2DD: out_word = 8'hFE;
		16'hA2DE: out_word = 8'hA5;
		16'hA2DF: out_word = 8'hC9;
		16'hA2E0: out_word = 8'h47;
		16'hA2E1: out_word = 8'hF6;
		16'hA2E2: out_word = 8'h20;
		16'hA2E3: out_word = 8'hFE;
		16'hA2E4: out_word = 8'h61;
		16'hA2E5: out_word = 8'h38;
		16'hA2E6: out_word = 8'h06;
		16'hA2E7: out_word = 8'hFE;
		16'hA2E8: out_word = 8'h7B;
		16'hA2E9: out_word = 8'h30;
		16'hA2EA: out_word = 8'h02;
		16'hA2EB: out_word = 8'hBF;
		16'hA2EC: out_word = 8'hC9;
		16'hA2ED: out_word = 8'h78;
		16'hA2EE: out_word = 8'hFE;
		16'hA2EF: out_word = 8'h2E;
		16'hA2F0: out_word = 8'hC8;
		16'hA2F1: out_word = 8'hCD;
		16'hA2F2: out_word = 8'h0A;
		16'hA2F3: out_word = 8'h23;
		16'hA2F4: out_word = 8'h20;
		16'hA2F5: out_word = 8'h11;
		16'hA2F6: out_word = 8'hE7;
		16'hA2F7: out_word = 8'hCD;
		16'hA2F8: out_word = 8'h0A;
		16'hA2F9: out_word = 8'h23;
		16'hA2FA: out_word = 8'h28;
		16'hA2FB: out_word = 8'hFA;
		16'hA2FC: out_word = 8'hFE;
		16'hA2FD: out_word = 8'h2E;
		16'hA2FE: out_word = 8'hC8;
		16'hA2FF: out_word = 8'hFE;
		16'hA300: out_word = 8'h45;
		16'hA301: out_word = 8'hC8;
		16'hA302: out_word = 8'hFE;
		16'hA303: out_word = 8'h65;
		16'hA304: out_word = 8'hC8;
		16'hA305: out_word = 8'h18;
		16'hA306: out_word = 8'hA4;
		16'hA307: out_word = 8'hF6;
		16'hA308: out_word = 8'hFF;
		16'hA309: out_word = 8'hC9;
		16'hA30A: out_word = 8'hFE;
		16'hA30B: out_word = 8'h30;
		16'hA30C: out_word = 8'h38;
		16'hA30D: out_word = 8'h06;
		16'hA30E: out_word = 8'hFE;
		16'hA30F: out_word = 8'h3A;
		16'hA310: out_word = 8'h30;
		16'hA311: out_word = 8'h02;
		16'hA312: out_word = 8'hBF;
		16'hA313: out_word = 8'hC9;
		16'hA314: out_word = 8'hFE;
		16'hA315: out_word = 8'h30;
		16'hA316: out_word = 8'hC9;
		16'hA317: out_word = 8'h06;
		16'hA318: out_word = 8'h00;
		16'hA319: out_word = 8'hDF;
		16'hA31A: out_word = 8'hC5;
		16'hA31B: out_word = 8'hEF;
		16'hA31C: out_word = 8'h8C;
		16'hA31D: out_word = 8'h1C;
		16'hA31E: out_word = 8'hC1;
		16'hA31F: out_word = 8'h04;
		16'hA320: out_word = 8'hFE;
		16'hA321: out_word = 8'h2C;
		16'hA322: out_word = 8'h20;
		16'hA323: out_word = 8'h03;
		16'hA324: out_word = 8'hE7;
		16'hA325: out_word = 8'h18;
		16'hA326: out_word = 8'hF3;
		16'hA327: out_word = 8'h78;
		16'hA328: out_word = 8'hFE;
		16'hA329: out_word = 8'h09;
		16'hA32A: out_word = 8'h38;
		16'hA32B: out_word = 8'h04;
		16'hA32C: out_word = 8'hCD;
		16'hA32D: out_word = 8'hAC;
		16'hA32E: out_word = 8'h05;
		16'hA32F: out_word = 8'h2B;
		16'hA330: out_word = 8'hCD;
		16'hA331: out_word = 8'hA1;
		16'hA332: out_word = 8'h18;
		16'hA333: out_word = 8'hC3;
		16'hA334: out_word = 8'h85;
		16'hA335: out_word = 8'h09;
		16'hA336: out_word = 8'h21;
		16'hA337: out_word = 8'hFF;
		16'hA338: out_word = 8'h5B;
		16'hA339: out_word = 8'h22;
		16'hA33A: out_word = 8'h81;
		16'hA33B: out_word = 8'h5B;
		16'hA33C: out_word = 8'hCD;
		16'hA33D: out_word = 8'h45;
		16'hA33E: out_word = 8'h1F;
		16'hA33F: out_word = 8'hC3;
		16'hA340: out_word = 8'hCB;
		16'hA341: out_word = 8'h25;
		16'hA342: out_word = 8'hA7;
		16'hA343: out_word = 8'hED;
		16'hA344: out_word = 8'h52;
		16'hA345: out_word = 8'h44;
		16'hA346: out_word = 8'h4D;
		16'hA347: out_word = 8'h19;
		16'hA348: out_word = 8'hEB;
		16'hA349: out_word = 8'hC9;
		16'hA34A: out_word = 8'h01;
		16'hA34B: out_word = 8'h01;
		16'hA34C: out_word = 8'h00;
		16'hA34D: out_word = 8'hE5;
		16'hA34E: out_word = 8'hD5;
		16'hA34F: out_word = 8'hCD;
		16'hA350: out_word = 8'h58;
		16'hA351: out_word = 8'h23;
		16'hA352: out_word = 8'hD1;
		16'hA353: out_word = 8'hE1;
		16'hA354: out_word = 8'hEF;
		16'hA355: out_word = 8'h55;
		16'hA356: out_word = 8'h16;
		16'hA357: out_word = 8'hC9;
		16'hA358: out_word = 8'h2A;
		16'hA359: out_word = 8'h65;
		16'hA35A: out_word = 8'h5C;
		16'hA35B: out_word = 8'h09;
		16'hA35C: out_word = 8'h38;
		16'hA35D: out_word = 8'h0A;
		16'hA35E: out_word = 8'hEB;
		16'hA35F: out_word = 8'h21;
		16'hA360: out_word = 8'h82;
		16'hA361: out_word = 8'h00;
		16'hA362: out_word = 8'h19;
		16'hA363: out_word = 8'h38;
		16'hA364: out_word = 8'h03;
		16'hA365: out_word = 8'hED;
		16'hA366: out_word = 8'h72;
		16'hA367: out_word = 8'hD8;
		16'hA368: out_word = 8'hFD;
		16'hA369: out_word = 8'h36;
		16'hA36A: out_word = 8'h00;
		16'hA36B: out_word = 8'h03;
		16'hA36C: out_word = 8'hC3;
		16'hA36D: out_word = 8'h21;
		16'hA36E: out_word = 8'h03;
		16'hA36F: out_word = 8'h87;
		16'hA370: out_word = 8'h87;
		16'hA371: out_word = 8'h6F;
		16'hA372: out_word = 8'h26;
		16'hA373: out_word = 8'h00;
		16'hA374: out_word = 8'h29;
		16'hA375: out_word = 8'h29;
		16'hA376: out_word = 8'h29;
		16'hA377: out_word = 8'hC9;
		16'hA378: out_word = 8'h21;
		16'hA379: out_word = 8'h00;
		16'hA37A: out_word = 8'h00;
		16'hA37B: out_word = 8'h39;
		16'hA37C: out_word = 8'hED;
		16'hA37D: out_word = 8'h5B;
		16'hA37E: out_word = 8'h65;
		16'hA37F: out_word = 8'h5C;
		16'hA380: out_word = 8'hB7;
		16'hA381: out_word = 8'hED;
		16'hA382: out_word = 8'h52;
		16'hA383: out_word = 8'hC9;
		16'hA384: out_word = 8'hFD;
		16'hA385: out_word = 8'hCB;
		16'hA386: out_word = 8'hC7;
		16'hA387: out_word = 8'h86;
		16'hA388: out_word = 8'hCD;
		16'hA389: out_word = 8'h6F;
		16'hA38A: out_word = 8'h23;
		16'hA38B: out_word = 8'hE5;
		16'hA38C: out_word = 8'hED;
		16'hA38D: out_word = 8'h5B;
		16'hA38E: out_word = 8'h24;
		16'hA38F: out_word = 8'hFF;
		16'hA390: out_word = 8'h19;
		16'hA391: out_word = 8'h54;
		16'hA392: out_word = 8'h5D;
		16'hA393: out_word = 8'hE3;
		16'hA394: out_word = 8'hE5;
		16'hA395: out_word = 8'hD5;
		16'hA396: out_word = 8'h11;
		16'hA397: out_word = 8'h00;
		16'hA398: out_word = 8'h58;
		16'hA399: out_word = 8'h19;
		16'hA39A: out_word = 8'hEB;
		16'hA39B: out_word = 8'hE1;
		16'hA39C: out_word = 8'h01;
		16'hA39D: out_word = 8'h20;
		16'hA39E: out_word = 8'h00;
		16'hA39F: out_word = 8'h3A;
		16'hA3A0: out_word = 8'h8F;
		16'hA3A1: out_word = 8'h5C;
		16'hA3A2: out_word = 8'hCD;
		16'hA3A3: out_word = 8'h9B;
		16'hA3A4: out_word = 8'h24;
		16'hA3A5: out_word = 8'hE1;
		16'hA3A6: out_word = 8'h7C;
		16'hA3A7: out_word = 8'h26;
		16'hA3A8: out_word = 8'h00;
		16'hA3A9: out_word = 8'h87;
		16'hA3AA: out_word = 8'h87;
		16'hA3AB: out_word = 8'h87;
		16'hA3AC: out_word = 8'hC6;
		16'hA3AD: out_word = 8'h40;
		16'hA3AE: out_word = 8'h57;
		16'hA3AF: out_word = 8'h5C;
		16'hA3B0: out_word = 8'h19;
		16'hA3B1: out_word = 8'hEB;
		16'hA3B2: out_word = 8'hE1;
		16'hA3B3: out_word = 8'h06;
		16'hA3B4: out_word = 8'h20;
		16'hA3B5: out_word = 8'hC3;
		16'hA3B6: out_word = 8'hE1;
		16'hA3B7: out_word = 8'h23;
		16'hA3B8: out_word = 8'h16;
		16'hA3B9: out_word = 8'hFF;
		16'hA3BA: out_word = 8'hCD;
		16'hA3BB: out_word = 8'h6F;
		16'hA3BC: out_word = 8'h23;
		16'hA3BD: out_word = 8'h7A;
		16'hA3BE: out_word = 8'hED;
		16'hA3BF: out_word = 8'h5B;
		16'hA3C0: out_word = 8'h24;
		16'hA3C1: out_word = 8'hFF;
		16'hA3C2: out_word = 8'h19;
		16'hA3C3: out_word = 8'h5D;
		16'hA3C4: out_word = 8'h54;
		16'hA3C5: out_word = 8'h13;
		16'hA3C6: out_word = 8'h77;
		16'hA3C7: out_word = 8'h0B;
		16'hA3C8: out_word = 8'hED;
		16'hA3C9: out_word = 8'hB0;
		16'hA3CA: out_word = 8'hC9;
		16'hA3CB: out_word = 8'hCD;
		16'hA3CC: out_word = 8'h88;
		16'hA3CD: out_word = 8'h24;
		16'hA3CE: out_word = 8'h11;
		16'hA3CF: out_word = 8'h00;
		16'hA3D0: out_word = 8'h40;
		16'hA3D1: out_word = 8'h2A;
		16'hA3D2: out_word = 8'h24;
		16'hA3D3: out_word = 8'hFF;
		16'hA3D4: out_word = 8'h43;
		16'hA3D5: out_word = 8'hCD;
		16'hA3D6: out_word = 8'hE1;
		16'hA3D7: out_word = 8'h23;
		16'hA3D8: out_word = 8'h16;
		16'hA3D9: out_word = 8'h48;
		16'hA3DA: out_word = 8'hCD;
		16'hA3DB: out_word = 8'hE1;
		16'hA3DC: out_word = 8'h23;
		16'hA3DD: out_word = 8'h16;
		16'hA3DE: out_word = 8'h50;
		16'hA3DF: out_word = 8'h06;
		16'hA3E0: out_word = 8'hC0;
		16'hA3E1: out_word = 8'h7E;
		16'hA3E2: out_word = 8'hE5;
		16'hA3E3: out_word = 8'hD5;
		16'hA3E4: out_word = 8'hFE;
		16'hA3E5: out_word = 8'hFE;
		16'hA3E6: out_word = 8'h38;
		16'hA3E7: out_word = 8'h04;
		16'hA3E8: out_word = 8'hD6;
		16'hA3E9: out_word = 8'hFE;
		16'hA3EA: out_word = 8'h18;
		16'hA3EB: out_word = 8'h36;
		16'hA3EC: out_word = 8'hFE;
		16'hA3ED: out_word = 8'h20;
		16'hA3EE: out_word = 8'h30;
		16'hA3EF: out_word = 8'h07;
		16'hA3F0: out_word = 8'h21;
		16'hA3F1: out_word = 8'h27;
		16'hA3F2: out_word = 8'h25;
		16'hA3F3: out_word = 8'hA7;
		16'hA3F4: out_word = 8'h08;
		16'hA3F5: out_word = 8'h18;
		16'hA3F6: out_word = 8'h34;
		16'hA3F7: out_word = 8'hFE;
		16'hA3F8: out_word = 8'h80;
		16'hA3F9: out_word = 8'h30;
		16'hA3FA: out_word = 8'h0E;
		16'hA3FB: out_word = 8'hCD;
		16'hA3FC: out_word = 8'h71;
		16'hA3FD: out_word = 8'h23;
		16'hA3FE: out_word = 8'hED;
		16'hA3FF: out_word = 8'h5B;
		16'hA400: out_word = 8'h36;
		16'hA401: out_word = 8'h5C;
		16'hA402: out_word = 8'h19;
		16'hA403: out_word = 8'hD1;
		16'hA404: out_word = 8'hCD;
		16'hA405: out_word = 8'h28;
		16'hA406: out_word = 8'hFF;
		16'hA407: out_word = 8'h18;
		16'hA408: out_word = 8'h47;
		16'hA409: out_word = 8'hFE;
		16'hA40A: out_word = 8'h90;
		16'hA40B: out_word = 8'h30;
		16'hA40C: out_word = 8'h04;
		16'hA40D: out_word = 8'hD6;
		16'hA40E: out_word = 8'h7F;
		16'hA40F: out_word = 8'h18;
		16'hA410: out_word = 8'h11;
		16'hA411: out_word = 8'hD6;
		16'hA412: out_word = 8'h90;
		16'hA413: out_word = 8'hCD;
		16'hA414: out_word = 8'h71;
		16'hA415: out_word = 8'h23;
		16'hA416: out_word = 8'hD1;
		16'hA417: out_word = 8'hCD;
		16'hA418: out_word = 8'h20;
		16'hA419: out_word = 8'h1F;
		16'hA41A: out_word = 8'hD5;
		16'hA41B: out_word = 8'hED;
		16'hA41C: out_word = 8'h5B;
		16'hA41D: out_word = 8'h7B;
		16'hA41E: out_word = 8'h5C;
		16'hA41F: out_word = 8'h37;
		16'hA420: out_word = 8'h18;
		16'hA421: out_word = 8'h07;
		16'hA422: out_word = 8'h11;
		16'hA423: out_word = 8'h2F;
		16'hA424: out_word = 8'h25;
		16'hA425: out_word = 8'hCD;
		16'hA426: out_word = 8'h71;
		16'hA427: out_word = 8'h23;
		16'hA428: out_word = 8'hA7;
		16'hA429: out_word = 8'h08;
		16'hA42A: out_word = 8'h19;
		16'hA42B: out_word = 8'hD1;
		16'hA42C: out_word = 8'h4A;
		16'hA42D: out_word = 8'h7E;
		16'hA42E: out_word = 8'h12;
		16'hA42F: out_word = 8'h23;
		16'hA430: out_word = 8'h14;
		16'hA431: out_word = 8'h7E;
		16'hA432: out_word = 8'h12;
		16'hA433: out_word = 8'h23;
		16'hA434: out_word = 8'h14;
		16'hA435: out_word = 8'h7E;
		16'hA436: out_word = 8'h12;
		16'hA437: out_word = 8'h23;
		16'hA438: out_word = 8'h14;
		16'hA439: out_word = 8'h7E;
		16'hA43A: out_word = 8'h12;
		16'hA43B: out_word = 8'h23;
		16'hA43C: out_word = 8'h14;
		16'hA43D: out_word = 8'h7E;
		16'hA43E: out_word = 8'h12;
		16'hA43F: out_word = 8'h23;
		16'hA440: out_word = 8'h14;
		16'hA441: out_word = 8'h7E;
		16'hA442: out_word = 8'h12;
		16'hA443: out_word = 8'h23;
		16'hA444: out_word = 8'h14;
		16'hA445: out_word = 8'h7E;
		16'hA446: out_word = 8'h12;
		16'hA447: out_word = 8'h23;
		16'hA448: out_word = 8'h14;
		16'hA449: out_word = 8'h7E;
		16'hA44A: out_word = 8'h12;
		16'hA44B: out_word = 8'h51;
		16'hA44C: out_word = 8'h08;
		16'hA44D: out_word = 8'hDC;
		16'hA44E: out_word = 8'h45;
		16'hA44F: out_word = 8'h1F;
		16'hA450: out_word = 8'hE1;
		16'hA451: out_word = 8'h23;
		16'hA452: out_word = 8'h13;
		16'hA453: out_word = 8'h10;
		16'hA454: out_word = 8'h8C;
		16'hA455: out_word = 8'hC9;
		16'hA456: out_word = 8'hC5;
		16'hA457: out_word = 8'hF3;
		16'hA458: out_word = 8'h01;
		16'hA459: out_word = 8'hFD;
		16'hA45A: out_word = 8'h7F;
		16'hA45B: out_word = 8'h3A;
		16'hA45C: out_word = 8'h5C;
		16'hA45D: out_word = 8'h5B;
		16'hA45E: out_word = 8'hEE;
		16'hA45F: out_word = 8'h10;
		16'hA460: out_word = 8'hED;
		16'hA461: out_word = 8'h79;
		16'hA462: out_word = 8'hFB;
		16'hA463: out_word = 8'h08;
		16'hA464: out_word = 8'h08;
		16'hA465: out_word = 8'hF3;
		16'hA466: out_word = 8'h0E;
		16'hA467: out_word = 8'hFD;
		16'hA468: out_word = 8'hEE;
		16'hA469: out_word = 8'h10;
		16'hA46A: out_word = 8'hED;
		16'hA46B: out_word = 8'h79;
		16'hA46C: out_word = 8'hFB;
		16'hA46D: out_word = 8'hC1;
		16'hA46E: out_word = 8'hC9;
		16'hA46F: out_word = 8'h21;
		16'hA470: out_word = 8'h56;
		16'hA471: out_word = 8'h24;
		16'hA472: out_word = 8'h11;
		16'hA473: out_word = 8'h28;
		16'hA474: out_word = 8'hFF;
		16'hA475: out_word = 8'h01;
		16'hA476: out_word = 8'h0E;
		16'hA477: out_word = 8'h00;
		16'hA478: out_word = 8'hED;
		16'hA479: out_word = 8'hB0;
		16'hA47A: out_word = 8'hE5;
		16'hA47B: out_word = 8'h21;
		16'hA47C: out_word = 8'h2C;
		16'hA47D: out_word = 8'h24;
		16'hA47E: out_word = 8'h0E;
		16'hA47F: out_word = 8'h20;
		16'hA480: out_word = 8'hED;
		16'hA481: out_word = 8'hB0;
		16'hA482: out_word = 8'hE1;
		16'hA483: out_word = 8'h0E;
		16'hA484: out_word = 8'h0B;
		16'hA485: out_word = 8'hED;
		16'hA486: out_word = 8'hB0;
		16'hA487: out_word = 8'hC9;
		16'hA488: out_word = 8'hFD;
		16'hA489: out_word = 8'hCB;
		16'hA48A: out_word = 8'hC7;
		16'hA48B: out_word = 8'h86;
		16'hA48C: out_word = 8'h11;
		16'hA48D: out_word = 8'h00;
		16'hA48E: out_word = 8'h58;
		16'hA48F: out_word = 8'h01;
		16'hA490: out_word = 8'hC0;
		16'hA491: out_word = 8'h02;
		16'hA492: out_word = 8'h2A;
		16'hA493: out_word = 8'h24;
		16'hA494: out_word = 8'hFF;
		16'hA495: out_word = 8'h3A;
		16'hA496: out_word = 8'h8D;
		16'hA497: out_word = 8'h5C;
		16'hA498: out_word = 8'h32;
		16'hA499: out_word = 8'h8F;
		16'hA49A: out_word = 8'h5C;
		16'hA49B: out_word = 8'h08;
		16'hA49C: out_word = 8'hC5;
		16'hA49D: out_word = 8'h7E;
		16'hA49E: out_word = 8'hFE;
		16'hA49F: out_word = 8'hFF;
		16'hA4A0: out_word = 8'h20;
		16'hA4A1: out_word = 8'h08;
		16'hA4A2: out_word = 8'h3A;
		16'hA4A3: out_word = 8'h8D;
		16'hA4A4: out_word = 8'h5C;
		16'hA4A5: out_word = 8'h12;
		16'hA4A6: out_word = 8'h23;
		16'hA4A7: out_word = 8'h13;
		16'hA4A8: out_word = 8'h18;
		16'hA4A9: out_word = 8'h5D;
		16'hA4AA: out_word = 8'h08;
		16'hA4AB: out_word = 8'h12;
		16'hA4AC: out_word = 8'h13;
		16'hA4AD: out_word = 8'h08;
		16'hA4AE: out_word = 8'h23;
		16'hA4AF: out_word = 8'hFE;
		16'hA4B0: out_word = 8'h15;
		16'hA4B1: out_word = 8'h30;
		16'hA4B2: out_word = 8'h54;
		16'hA4B3: out_word = 8'hFE;
		16'hA4B4: out_word = 8'h10;
		16'hA4B5: out_word = 8'h38;
		16'hA4B6: out_word = 8'h50;
		16'hA4B7: out_word = 8'h2B;
		16'hA4B8: out_word = 8'h20;
		16'hA4B9: out_word = 8'h08;
		16'hA4BA: out_word = 8'h23;
		16'hA4BB: out_word = 8'h7E;
		16'hA4BC: out_word = 8'h4F;
		16'hA4BD: out_word = 8'h08;
		16'hA4BE: out_word = 8'hE6;
		16'hA4BF: out_word = 8'hF8;
		16'hA4C0: out_word = 8'h18;
		16'hA4C1: out_word = 8'h43;
		16'hA4C2: out_word = 8'hFE;
		16'hA4C3: out_word = 8'h11;
		16'hA4C4: out_word = 8'h20;
		16'hA4C5: out_word = 8'h0B;
		16'hA4C6: out_word = 8'h23;
		16'hA4C7: out_word = 8'h7E;
		16'hA4C8: out_word = 8'h87;
		16'hA4C9: out_word = 8'h87;
		16'hA4CA: out_word = 8'h87;
		16'hA4CB: out_word = 8'h4F;
		16'hA4CC: out_word = 8'h08;
		16'hA4CD: out_word = 8'hE6;
		16'hA4CE: out_word = 8'hC7;
		16'hA4CF: out_word = 8'h18;
		16'hA4D0: out_word = 8'h34;
		16'hA4D1: out_word = 8'hFE;
		16'hA4D2: out_word = 8'h12;
		16'hA4D3: out_word = 8'h20;
		16'hA4D4: out_word = 8'h09;
		16'hA4D5: out_word = 8'h23;
		16'hA4D6: out_word = 8'h7E;
		16'hA4D7: out_word = 8'h0F;
		16'hA4D8: out_word = 8'h4F;
		16'hA4D9: out_word = 8'h08;
		16'hA4DA: out_word = 8'hE6;
		16'hA4DB: out_word = 8'h7F;
		16'hA4DC: out_word = 8'h18;
		16'hA4DD: out_word = 8'h27;
		16'hA4DE: out_word = 8'hFE;
		16'hA4DF: out_word = 8'h13;
		16'hA4E0: out_word = 8'h20;
		16'hA4E1: out_word = 8'h0A;
		16'hA4E2: out_word = 8'h23;
		16'hA4E3: out_word = 8'h7E;
		16'hA4E4: out_word = 8'h0F;
		16'hA4E5: out_word = 8'h0F;
		16'hA4E6: out_word = 8'h4F;
		16'hA4E7: out_word = 8'h08;
		16'hA4E8: out_word = 8'hE6;
		16'hA4E9: out_word = 8'hBF;
		16'hA4EA: out_word = 8'h18;
		16'hA4EB: out_word = 8'h19;
		16'hA4EC: out_word = 8'hFE;
		16'hA4ED: out_word = 8'h14;
		16'hA4EE: out_word = 8'h23;
		16'hA4EF: out_word = 8'h20;
		16'hA4F0: out_word = 8'h16;
		16'hA4F1: out_word = 8'h4E;
		16'hA4F2: out_word = 8'h3A;
		16'hA4F3: out_word = 8'h01;
		16'hA4F4: out_word = 8'h5C;
		16'hA4F5: out_word = 8'hA9;
		16'hA4F6: out_word = 8'h1F;
		16'hA4F7: out_word = 8'h30;
		16'hA4F8: out_word = 8'h0E;
		16'hA4F9: out_word = 8'h3E;
		16'hA4FA: out_word = 8'h01;
		16'hA4FB: out_word = 8'hFD;
		16'hA4FC: out_word = 8'hAE;
		16'hA4FD: out_word = 8'hC7;
		16'hA4FE: out_word = 8'h32;
		16'hA4FF: out_word = 8'h01;
		16'hA500: out_word = 8'h5C;
		16'hA501: out_word = 8'h08;
		16'hA502: out_word = 8'hCD;
		16'hA503: out_word = 8'h13;
		16'hA504: out_word = 8'h25;
		16'hA505: out_word = 8'hB1;
		16'hA506: out_word = 8'h08;
		16'hA507: out_word = 8'hC1;
		16'hA508: out_word = 8'h0B;
		16'hA509: out_word = 8'h78;
		16'hA50A: out_word = 8'hB1;
		16'hA50B: out_word = 8'hC2;
		16'hA50C: out_word = 8'h9C;
		16'hA50D: out_word = 8'h24;
		16'hA50E: out_word = 8'h08;
		16'hA50F: out_word = 8'h32;
		16'hA510: out_word = 8'h8F;
		16'hA511: out_word = 8'h5C;
		16'hA512: out_word = 8'hC9;
		16'hA513: out_word = 8'h47;
		16'hA514: out_word = 8'hE6;
		16'hA515: out_word = 8'hC0;
		16'hA516: out_word = 8'h4F;
		16'hA517: out_word = 8'h78;
		16'hA518: out_word = 8'h87;
		16'hA519: out_word = 8'h87;
		16'hA51A: out_word = 8'h87;
		16'hA51B: out_word = 8'hE6;
		16'hA51C: out_word = 8'h38;
		16'hA51D: out_word = 8'hB1;
		16'hA51E: out_word = 8'h4F;
		16'hA51F: out_word = 8'h78;
		16'hA520: out_word = 8'h1F;
		16'hA521: out_word = 8'h1F;
		16'hA522: out_word = 8'h1F;
		16'hA523: out_word = 8'hE6;
		16'hA524: out_word = 8'h07;
		16'hA525: out_word = 8'hB1;
		16'hA526: out_word = 8'hC9;
		16'hA527: out_word = 8'h00;
		16'hA528: out_word = 8'h3C;
		16'hA529: out_word = 8'h62;
		16'hA52A: out_word = 8'h60;
		16'hA52B: out_word = 8'h6E;
		16'hA52C: out_word = 8'h62;
		16'hA52D: out_word = 8'h3E;
		16'hA52E: out_word = 8'h00;
		16'hA52F: out_word = 8'h00;
		16'hA530: out_word = 8'h6C;
		16'hA531: out_word = 8'h10;
		16'hA532: out_word = 8'h54;
		16'hA533: out_word = 8'hBA;
		16'hA534: out_word = 8'h38;
		16'hA535: out_word = 8'h54;
		16'hA536: out_word = 8'h82;
		16'hA537: out_word = 8'h15;
		16'hA538: out_word = 8'h0B;
		16'hA539: out_word = 8'h94;
		16'hA53A: out_word = 8'h2A;
		16'hA53B: out_word = 8'h0A;
		16'hA53C: out_word = 8'hB5;
		16'hA53D: out_word = 8'h2A;
		16'hA53E: out_word = 8'h08;
		16'hA53F: out_word = 8'hD7;
		16'hA540: out_word = 8'h2A;
		16'hA541: out_word = 8'h09;
		16'hA542: out_word = 8'hE3;
		16'hA543: out_word = 8'h2A;
		16'hA544: out_word = 8'hAD;
		16'hA545: out_word = 8'h4F;
		16'hA546: out_word = 8'h2A;
		16'hA547: out_word = 8'hAC;
		16'hA548: out_word = 8'h25;
		16'hA549: out_word = 8'h2A;
		16'hA54A: out_word = 8'hAF;
		16'hA54B: out_word = 8'hD4;
		16'hA54C: out_word = 8'h29;
		16'hA54D: out_word = 8'hAE;
		16'hA54E: out_word = 8'hE1;
		16'hA54F: out_word = 8'h29;
		16'hA550: out_word = 8'hA6;
		16'hA551: out_word = 8'h83;
		16'hA552: out_word = 8'h29;
		16'hA553: out_word = 8'hA5;
		16'hA554: out_word = 8'hAB;
		16'hA555: out_word = 8'h29;
		16'hA556: out_word = 8'hA8;
		16'hA557: out_word = 8'h87;
		16'hA558: out_word = 8'h2A;
		16'hA559: out_word = 8'hA7;
		16'hA55A: out_word = 8'h7A;
		16'hA55B: out_word = 8'h2A;
		16'hA55C: out_word = 8'hAA;
		16'hA55D: out_word = 8'h1B;
		16'hA55E: out_word = 8'h29;
		16'hA55F: out_word = 8'h0C;
		16'hA560: out_word = 8'h2B;
		16'hA561: out_word = 8'h29;
		16'hA562: out_word = 8'hB3;
		16'hA563: out_word = 8'h17;
		16'hA564: out_word = 8'h30;
		16'hA565: out_word = 8'hB4;
		16'hA566: out_word = 8'hBC;
		16'hA567: out_word = 8'h2F;
		16'hA568: out_word = 8'hB0;
		16'hA569: out_word = 8'h72;
		16'hA56A: out_word = 8'h30;
		16'hA56B: out_word = 8'hB1;
		16'hA56C: out_word = 8'h3E;
		16'hA56D: out_word = 8'h30;
		16'hA56E: out_word = 8'h0D;
		16'hA56F: out_word = 8'h44;
		16'hA570: out_word = 8'h29;
		16'hA571: out_word = 8'hA9;
		16'hA572: out_word = 8'h9B;
		16'hA573: out_word = 8'h26;
		16'hA574: out_word = 8'h07;
		16'hA575: out_word = 8'h04;
		16'hA576: out_word = 8'h27;
		16'hA577: out_word = 8'h04;
		16'hA578: out_word = 8'h0B;
		16'hA579: out_word = 8'h2E;
		16'hA57A: out_word = 8'h27;
		16'hA57B: out_word = 8'h0A;
		16'hA57C: out_word = 8'h31;
		16'hA57D: out_word = 8'h27;
		16'hA57E: out_word = 8'h07;
		16'hA57F: out_word = 8'h17;
		16'hA580: out_word = 8'h27;
		16'hA581: out_word = 8'h0D;
		16'hA582: out_word = 8'h17;
		16'hA583: out_word = 8'h27;
		16'hA584: out_word = 8'hCD;
		16'hA585: out_word = 8'hBE;
		16'hA586: out_word = 8'h28;
		16'hA587: out_word = 8'h21;
		16'hA588: out_word = 8'h00;
		16'hA589: out_word = 8'h00;
		16'hA58A: out_word = 8'h22;
		16'hA58B: out_word = 8'h9A;
		16'hA58C: out_word = 8'hFC;
		16'hA58D: out_word = 8'h3E;
		16'hA58E: out_word = 8'h82;
		16'hA58F: out_word = 8'h32;
		16'hA590: out_word = 8'h0D;
		16'hA591: out_word = 8'hEC;
		16'hA592: out_word = 8'h21;
		16'hA593: out_word = 8'h00;
		16'hA594: out_word = 8'h00;
		16'hA595: out_word = 8'h22;
		16'hA596: out_word = 8'h49;
		16'hA597: out_word = 8'h5C;
		16'hA598: out_word = 8'hCD;
		16'hA599: out_word = 8'hBC;
		16'hA59A: out_word = 8'h35;
		16'hA59B: out_word = 8'hCD;
		16'hA59C: out_word = 8'h5E;
		16'hA59D: out_word = 8'h36;
		16'hA59E: out_word = 8'hC9;
		16'hA59F: out_word = 8'h21;
		16'hA5A0: out_word = 8'hFF;
		16'hA5A1: out_word = 8'h5B;
		16'hA5A2: out_word = 8'h22;
		16'hA5A3: out_word = 8'h81;
		16'hA5A4: out_word = 8'h5B;
		16'hA5A5: out_word = 8'hCD;
		16'hA5A6: out_word = 8'h45;
		16'hA5A7: out_word = 8'h1F;
		16'hA5A8: out_word = 8'h3E;
		16'hA5A9: out_word = 8'h02;
		16'hA5AA: out_word = 8'hEF;
		16'hA5AB: out_word = 8'h01;
		16'hA5AC: out_word = 8'h16;
		16'hA5AD: out_word = 8'h21;
		16'hA5AE: out_word = 8'h44;
		16'hA5AF: out_word = 8'h27;
		16'hA5B0: out_word = 8'h22;
		16'hA5B1: out_word = 8'hEA;
		16'hA5B2: out_word = 8'hF6;
		16'hA5B3: out_word = 8'h21;
		16'hA5B4: out_word = 8'h54;
		16'hA5B5: out_word = 8'h27;
		16'hA5B6: out_word = 8'h22;
		16'hA5B7: out_word = 8'hEC;
		16'hA5B8: out_word = 8'hF6;
		16'hA5B9: out_word = 8'hE5;
		16'hA5BA: out_word = 8'h21;
		16'hA5BB: out_word = 8'h0D;
		16'hA5BC: out_word = 8'hEC;
		16'hA5BD: out_word = 8'hCB;
		16'hA5BE: out_word = 8'hCE;
		16'hA5BF: out_word = 8'hCB;
		16'hA5C0: out_word = 8'hA6;
		16'hA5C1: out_word = 8'h2B;
		16'hA5C2: out_word = 8'h36;
		16'hA5C3: out_word = 8'h00;
		16'hA5C4: out_word = 8'hE1;
		16'hA5C5: out_word = 8'hCD;
		16'hA5C6: out_word = 8'hA8;
		16'hA5C7: out_word = 8'h36;
		16'hA5C8: out_word = 8'hC3;
		16'hA5C9: out_word = 8'h53;
		16'hA5CA: out_word = 8'h26;
		16'hA5CB: out_word = 8'hDD;
		16'hA5CC: out_word = 8'h21;
		16'hA5CD: out_word = 8'h6C;
		16'hA5CE: out_word = 8'hFD;
		16'hA5CF: out_word = 8'h21;
		16'hA5D0: out_word = 8'hFF;
		16'hA5D1: out_word = 8'h5B;
		16'hA5D2: out_word = 8'h22;
		16'hA5D3: out_word = 8'h81;
		16'hA5D4: out_word = 8'h5B;
		16'hA5D5: out_word = 8'hCD;
		16'hA5D6: out_word = 8'h45;
		16'hA5D7: out_word = 8'h1F;
		16'hA5D8: out_word = 8'h3E;
		16'hA5D9: out_word = 8'h02;
		16'hA5DA: out_word = 8'hEF;
		16'hA5DB: out_word = 8'h01;
		16'hA5DC: out_word = 8'h16;
		16'hA5DD: out_word = 8'hCD;
		16'hA5DE: out_word = 8'h68;
		16'hA5DF: out_word = 8'h36;
		16'hA5E0: out_word = 8'h21;
		16'hA5E1: out_word = 8'h3B;
		16'hA5E2: out_word = 8'h5C;
		16'hA5E3: out_word = 8'hCB;
		16'hA5E4: out_word = 8'h6E;
		16'hA5E5: out_word = 8'h28;
		16'hA5E6: out_word = 8'hFC;
		16'hA5E7: out_word = 8'h21;
		16'hA5E8: out_word = 8'h0D;
		16'hA5E9: out_word = 8'hEC;
		16'hA5EA: out_word = 8'hCB;
		16'hA5EB: out_word = 8'h9E;
		16'hA5EC: out_word = 8'hCB;
		16'hA5ED: out_word = 8'h76;
		16'hA5EE: out_word = 8'h20;
		16'hA5EF: out_word = 8'h14;
		16'hA5F0: out_word = 8'h3A;
		16'hA5F1: out_word = 8'h0E;
		16'hA5F2: out_word = 8'hEC;
		16'hA5F3: out_word = 8'hFE;
		16'hA5F4: out_word = 8'h04;
		16'hA5F5: out_word = 8'h28;
		16'hA5F6: out_word = 8'h0A;
		16'hA5F7: out_word = 8'hFE;
		16'hA5F8: out_word = 8'h00;
		16'hA5F9: out_word = 8'hC2;
		16'hA5FA: out_word = 8'hC7;
		16'hA5FB: out_word = 8'h28;
		16'hA5FC: out_word = 8'hCD;
		16'hA5FD: out_word = 8'h48;
		16'hA5FE: out_word = 8'h38;
		16'hA5FF: out_word = 8'h18;
		16'hA600: out_word = 8'h03;
		16'hA601: out_word = 8'hCD;
		16'hA602: out_word = 8'h4D;
		16'hA603: out_word = 8'h38;
		16'hA604: out_word = 8'hCD;
		16'hA605: out_word = 8'hD6;
		16'hA606: out_word = 8'h30;
		16'hA607: out_word = 8'hCD;
		16'hA608: out_word = 8'h22;
		16'hA609: out_word = 8'h32;
		16'hA60A: out_word = 8'h3A;
		16'hA60B: out_word = 8'h0E;
		16'hA60C: out_word = 8'hEC;
		16'hA60D: out_word = 8'hFE;
		16'hA60E: out_word = 8'h04;
		16'hA60F: out_word = 8'h28;
		16'hA610: out_word = 8'h42;
		16'hA611: out_word = 8'h2A;
		16'hA612: out_word = 8'h49;
		16'hA613: out_word = 8'h5C;
		16'hA614: out_word = 8'h7C;
		16'hA615: out_word = 8'hB5;
		16'hA616: out_word = 8'h20;
		16'hA617: out_word = 8'h15;
		16'hA618: out_word = 8'h2A;
		16'hA619: out_word = 8'h53;
		16'hA61A: out_word = 8'h5C;
		16'hA61B: out_word = 8'hED;
		16'hA61C: out_word = 8'h4B;
		16'hA61D: out_word = 8'h4B;
		16'hA61E: out_word = 8'h5C;
		16'hA61F: out_word = 8'hA7;
		16'hA620: out_word = 8'hED;
		16'hA621: out_word = 8'h42;
		16'hA622: out_word = 8'h20;
		16'hA623: out_word = 8'h06;
		16'hA624: out_word = 8'h21;
		16'hA625: out_word = 8'h00;
		16'hA626: out_word = 8'h00;
		16'hA627: out_word = 8'h22;
		16'hA628: out_word = 8'h08;
		16'hA629: out_word = 8'hEC;
		16'hA62A: out_word = 8'h2A;
		16'hA62B: out_word = 8'h08;
		16'hA62C: out_word = 8'hEC;
		16'hA62D: out_word = 8'hCD;
		16'hA62E: out_word = 8'h20;
		16'hA62F: out_word = 8'h1F;
		16'hA630: out_word = 8'hEF;
		16'hA631: out_word = 8'h6E;
		16'hA632: out_word = 8'h19;
		16'hA633: out_word = 8'hEF;
		16'hA634: out_word = 8'h95;
		16'hA635: out_word = 8'h16;
		16'hA636: out_word = 8'hCD;
		16'hA637: out_word = 8'h45;
		16'hA638: out_word = 8'h1F;
		16'hA639: out_word = 8'hED;
		16'hA63A: out_word = 8'h53;
		16'hA63B: out_word = 8'h49;
		16'hA63C: out_word = 8'h5C;
		16'hA63D: out_word = 8'h21;
		16'hA63E: out_word = 8'h0D;
		16'hA63F: out_word = 8'hEC;
		16'hA640: out_word = 8'hCB;
		16'hA641: out_word = 8'h6E;
		16'hA642: out_word = 8'h20;
		16'hA643: out_word = 8'h0F;
		16'hA644: out_word = 8'h21;
		16'hA645: out_word = 8'h00;
		16'hA646: out_word = 8'h00;
		16'hA647: out_word = 8'h22;
		16'hA648: out_word = 8'h06;
		16'hA649: out_word = 8'hEC;
		16'hA64A: out_word = 8'hCD;
		16'hA64B: out_word = 8'h2F;
		16'hA64C: out_word = 8'h15;
		16'hA64D: out_word = 8'hCD;
		16'hA64E: out_word = 8'hF2;
		16'hA64F: out_word = 8'h29;
		16'hA650: out_word = 8'hCD;
		16'hA651: out_word = 8'h44;
		16'hA652: out_word = 8'h29;
		16'hA653: out_word = 8'h31;
		16'hA654: out_word = 8'hFF;
		16'hA655: out_word = 8'h5B;
		16'hA656: out_word = 8'hCD;
		16'hA657: out_word = 8'h68;
		16'hA658: out_word = 8'h36;
		16'hA659: out_word = 8'hCD;
		16'hA65A: out_word = 8'h7F;
		16'hA65B: out_word = 8'h36;
		16'hA65C: out_word = 8'hF5;
		16'hA65D: out_word = 8'h3A;
		16'hA65E: out_word = 8'h39;
		16'hA65F: out_word = 8'h5C;
		16'hA660: out_word = 8'hCD;
		16'hA661: out_word = 8'hEC;
		16'hA662: out_word = 8'h26;
		16'hA663: out_word = 8'hF1;
		16'hA664: out_word = 8'hCD;
		16'hA665: out_word = 8'h69;
		16'hA666: out_word = 8'h26;
		16'hA667: out_word = 8'h18;
		16'hA668: out_word = 8'hEA;
		16'hA669: out_word = 8'h21;
		16'hA66A: out_word = 8'h0D;
		16'hA66B: out_word = 8'hEC;
		16'hA66C: out_word = 8'hCB;
		16'hA66D: out_word = 8'h4E;
		16'hA66E: out_word = 8'hF5;
		16'hA66F: out_word = 8'h21;
		16'hA670: out_word = 8'h77;
		16'hA671: out_word = 8'h25;
		16'hA672: out_word = 8'h20;
		16'hA673: out_word = 8'h03;
		16'hA674: out_word = 8'h21;
		16'hA675: out_word = 8'h37;
		16'hA676: out_word = 8'h25;
		16'hA677: out_word = 8'hCD;
		16'hA678: out_word = 8'hCE;
		16'hA679: out_word = 8'h3F;
		16'hA67A: out_word = 8'h20;
		16'hA67B: out_word = 8'h05;
		16'hA67C: out_word = 8'hD4;
		16'hA67D: out_word = 8'hE7;
		16'hA67E: out_word = 8'h26;
		16'hA67F: out_word = 8'hF1;
		16'hA680: out_word = 8'hC9;
		16'hA681: out_word = 8'hF1;
		16'hA682: out_word = 8'h28;
		16'hA683: out_word = 8'h05;
		16'hA684: out_word = 8'hAF;
		16'hA685: out_word = 8'h32;
		16'hA686: out_word = 8'h41;
		16'hA687: out_word = 8'h5C;
		16'hA688: out_word = 8'hC9;
		16'hA689: out_word = 8'h21;
		16'hA68A: out_word = 8'h0D;
		16'hA68B: out_word = 8'hEC;
		16'hA68C: out_word = 8'hCB;
		16'hA68D: out_word = 8'h46;
		16'hA68E: out_word = 8'h28;
		16'hA68F: out_word = 8'h04;
		16'hA690: out_word = 8'hCD;
		16'hA691: out_word = 8'hE7;
		16'hA692: out_word = 8'h26;
		16'hA693: out_word = 8'hC9;
		16'hA694: out_word = 8'hFE;
		16'hA695: out_word = 8'hA3;
		16'hA696: out_word = 8'h30;
		16'hA697: out_word = 8'hBB;
		16'hA698: out_word = 8'hC3;
		16'hA699: out_word = 8'hF1;
		16'hA69A: out_word = 8'h28;
		16'hA69B: out_word = 8'h3A;
		16'hA69C: out_word = 8'h0E;
		16'hA69D: out_word = 8'hEC;
		16'hA69E: out_word = 8'hFE;
		16'hA69F: out_word = 8'h04;
		16'hA6A0: out_word = 8'hC8;
		16'hA6A1: out_word = 8'hCD;
		16'hA6A2: out_word = 8'h30;
		16'hA6A3: out_word = 8'h16;
		16'hA6A4: out_word = 8'h21;
		16'hA6A5: out_word = 8'h0D;
		16'hA6A6: out_word = 8'hEC;
		16'hA6A7: out_word = 8'hCB;
		16'hA6A8: out_word = 8'h9E;
		16'hA6A9: out_word = 8'h7E;
		16'hA6AA: out_word = 8'hEE;
		16'hA6AB: out_word = 8'h40;
		16'hA6AC: out_word = 8'h77;
		16'hA6AD: out_word = 8'hE6;
		16'hA6AE: out_word = 8'h40;
		16'hA6AF: out_word = 8'h28;
		16'hA6B0: out_word = 8'h05;
		16'hA6B1: out_word = 8'hCD;
		16'hA6B2: out_word = 8'hBB;
		16'hA6B3: out_word = 8'h26;
		16'hA6B4: out_word = 8'h18;
		16'hA6B5: out_word = 8'h03;
		16'hA6B6: out_word = 8'hCD;
		16'hA6B7: out_word = 8'hCE;
		16'hA6B8: out_word = 8'h26;
		16'hA6B9: out_word = 8'h37;
		16'hA6BA: out_word = 8'hC9;
		16'hA6BB: out_word = 8'hCD;
		16'hA6BC: out_word = 8'h81;
		16'hA6BD: out_word = 8'h38;
		16'hA6BE: out_word = 8'h21;
		16'hA6BF: out_word = 8'h0D;
		16'hA6C0: out_word = 8'hEC;
		16'hA6C1: out_word = 8'hCB;
		16'hA6C2: out_word = 8'hF6;
		16'hA6C3: out_word = 8'hCD;
		16'hA6C4: out_word = 8'h2D;
		16'hA6C5: out_word = 8'h2E;
		16'hA6C6: out_word = 8'hCD;
		16'hA6C7: out_word = 8'h88;
		16'hA6C8: out_word = 8'h3A;
		16'hA6C9: out_word = 8'hCD;
		16'hA6CA: out_word = 8'hDF;
		16'hA6CB: out_word = 8'h28;
		16'hA6CC: out_word = 8'h18;
		16'hA6CD: out_word = 8'h0B;
		16'hA6CE: out_word = 8'h21;
		16'hA6CF: out_word = 8'h0D;
		16'hA6D0: out_word = 8'hEC;
		16'hA6D1: out_word = 8'hCB;
		16'hA6D2: out_word = 8'hB6;
		16'hA6D3: out_word = 8'hCD;
		16'hA6D4: out_word = 8'hBE;
		16'hA6D5: out_word = 8'h28;
		16'hA6D6: out_word = 8'hCD;
		16'hA6D7: out_word = 8'h48;
		16'hA6D8: out_word = 8'h38;
		16'hA6D9: out_word = 8'h2A;
		16'hA6DA: out_word = 8'h9A;
		16'hA6DB: out_word = 8'hFC;
		16'hA6DC: out_word = 8'h7C;
		16'hA6DD: out_word = 8'hB5;
		16'hA6DE: out_word = 8'hC4;
		16'hA6DF: out_word = 8'h4A;
		16'hA6E0: out_word = 8'h33;
		16'hA6E1: out_word = 8'hCD;
		16'hA6E2: out_word = 8'h2F;
		16'hA6E3: out_word = 8'h15;
		16'hA6E4: out_word = 8'hC3;
		16'hA6E5: out_word = 8'hF2;
		16'hA6E6: out_word = 8'h29;
		16'hA6E7: out_word = 8'h3A;
		16'hA6E8: out_word = 8'h38;
		16'hA6E9: out_word = 8'h5C;
		16'hA6EA: out_word = 8'hCB;
		16'hA6EB: out_word = 8'h3F;
		16'hA6EC: out_word = 8'hDD;
		16'hA6ED: out_word = 8'hE5;
		16'hA6EE: out_word = 8'h16;
		16'hA6EF: out_word = 8'h00;
		16'hA6F0: out_word = 8'h5F;
		16'hA6F1: out_word = 8'h21;
		16'hA6F2: out_word = 8'h80;
		16'hA6F3: out_word = 8'h0C;
		16'hA6F4: out_word = 8'hEF;
		16'hA6F5: out_word = 8'hB5;
		16'hA6F6: out_word = 8'h03;
		16'hA6F7: out_word = 8'hDD;
		16'hA6F8: out_word = 8'hE1;
		16'hA6F9: out_word = 8'hC9;
		16'hA6FA: out_word = 8'hDD;
		16'hA6FB: out_word = 8'hE5;
		16'hA6FC: out_word = 8'h11;
		16'hA6FD: out_word = 8'h30;
		16'hA6FE: out_word = 8'h00;
		16'hA6FF: out_word = 8'h21;
		16'hA700: out_word = 8'h00;
		16'hA701: out_word = 8'h03;
		16'hA702: out_word = 8'h18;
		16'hA703: out_word = 8'hF0;
		16'hA704: out_word = 8'hCD;
		16'hA705: out_word = 8'hEC;
		16'hA706: out_word = 8'h29;
		16'hA707: out_word = 8'h21;
		16'hA708: out_word = 8'h0D;
		16'hA709: out_word = 8'hEC;
		16'hA70A: out_word = 8'hCB;
		16'hA70B: out_word = 8'hCE;
		16'hA70C: out_word = 8'h2B;
		16'hA70D: out_word = 8'h36;
		16'hA70E: out_word = 8'h00;
		16'hA70F: out_word = 8'h2A;
		16'hA710: out_word = 8'hEC;
		16'hA711: out_word = 8'hF6;
		16'hA712: out_word = 8'hCD;
		16'hA713: out_word = 8'hA8;
		16'hA714: out_word = 8'h36;
		16'hA715: out_word = 8'h37;
		16'hA716: out_word = 8'hC9;
		16'hA717: out_word = 8'h21;
		16'hA718: out_word = 8'h0D;
		16'hA719: out_word = 8'hEC;
		16'hA71A: out_word = 8'hCB;
		16'hA71B: out_word = 8'h8E;
		16'hA71C: out_word = 8'h2B;
		16'hA71D: out_word = 8'h7E;
		16'hA71E: out_word = 8'h2A;
		16'hA71F: out_word = 8'hEA;
		16'hA720: out_word = 8'hF6;
		16'hA721: out_word = 8'hE5;
		16'hA722: out_word = 8'hF5;
		16'hA723: out_word = 8'hCD;
		16'hA724: out_word = 8'h3E;
		16'hA725: out_word = 8'h37;
		16'hA726: out_word = 8'hF1;
		16'hA727: out_word = 8'hE1;
		16'hA728: out_word = 8'hCD;
		16'hA729: out_word = 8'hCE;
		16'hA72A: out_word = 8'h3F;
		16'hA72B: out_word = 8'hC3;
		16'hA72C: out_word = 8'hF2;
		16'hA72D: out_word = 8'h29;
		16'hA72E: out_word = 8'h37;
		16'hA72F: out_word = 8'h18;
		16'hA730: out_word = 8'h01;
		16'hA731: out_word = 8'hA7;
		16'hA732: out_word = 8'h21;
		16'hA733: out_word = 8'h0C;
		16'hA734: out_word = 8'hEC;
		16'hA735: out_word = 8'h7E;
		16'hA736: out_word = 8'hE5;
		16'hA737: out_word = 8'h2A;
		16'hA738: out_word = 8'hEC;
		16'hA739: out_word = 8'hF6;
		16'hA73A: out_word = 8'hDC;
		16'hA73B: out_word = 8'hA7;
		16'hA73C: out_word = 8'h37;
		16'hA73D: out_word = 8'hD4;
		16'hA73E: out_word = 8'hB6;
		16'hA73F: out_word = 8'h37;
		16'hA740: out_word = 8'hE1;
		16'hA741: out_word = 8'h77;
		16'hA742: out_word = 8'h37;
		16'hA743: out_word = 8'hC9;
		16'hA744: out_word = 8'h05;
		16'hA745: out_word = 8'h00;
		16'hA746: out_word = 8'h31;
		16'hA747: out_word = 8'h28;
		16'hA748: out_word = 8'h01;
		16'hA749: out_word = 8'h6C;
		16'hA74A: out_word = 8'h28;
		16'hA74B: out_word = 8'h02;
		16'hA74C: out_word = 8'h85;
		16'hA74D: out_word = 8'h28;
		16'hA74E: out_word = 8'h03;
		16'hA74F: out_word = 8'h47;
		16'hA750: out_word = 8'h1B;
		16'hA751: out_word = 8'h04;
		16'hA752: out_word = 8'h16;
		16'hA753: out_word = 8'h28;
		16'hA754: out_word = 8'h06;
		16'hA755: out_word = 8'h31;
		16'hA756: out_word = 8'h32;
		16'hA757: out_word = 8'h38;
		16'hA758: out_word = 8'h20;
		16'hA759: out_word = 8'h20;
		16'hA75A: out_word = 8'h20;
		16'hA75B: out_word = 8'h20;
		16'hA75C: out_word = 8'h20;
		16'hA75D: out_word = 8'hFF;
		16'hA75E: out_word = 8'h54;
		16'hA75F: out_word = 8'h61;
		16'hA760: out_word = 8'h70;
		16'hA761: out_word = 8'h65;
		16'hA762: out_word = 8'h20;
		16'hA763: out_word = 8'h4C;
		16'hA764: out_word = 8'h6F;
		16'hA765: out_word = 8'h61;
		16'hA766: out_word = 8'h64;
		16'hA767: out_word = 8'h65;
		16'hA768: out_word = 8'hF2;
		16'hA769: out_word = 8'h31;
		16'hA76A: out_word = 8'h32;
		16'hA76B: out_word = 8'h38;
		16'hA76C: out_word = 8'h20;
		16'hA76D: out_word = 8'h42;
		16'hA76E: out_word = 8'h41;
		16'hA76F: out_word = 8'h53;
		16'hA770: out_word = 8'h49;
		16'hA771: out_word = 8'hC3;
		16'hA772: out_word = 8'h43;
		16'hA773: out_word = 8'h61;
		16'hA774: out_word = 8'h6C;
		16'hA775: out_word = 8'h63;
		16'hA776: out_word = 8'h75;
		16'hA777: out_word = 8'h6C;
		16'hA778: out_word = 8'h61;
		16'hA779: out_word = 8'h74;
		16'hA77A: out_word = 8'h6F;
		16'hA77B: out_word = 8'hF2;
		16'hA77C: out_word = 8'h34;
		16'hA77D: out_word = 8'h38;
		16'hA77E: out_word = 8'h20;
		16'hA77F: out_word = 8'h42;
		16'hA780: out_word = 8'h41;
		16'hA781: out_word = 8'h53;
		16'hA782: out_word = 8'h49;
		16'hA783: out_word = 8'hC3;
		16'hA784: out_word = 8'h54;
		16'hA785: out_word = 8'h52;
		16'hA786: out_word = 8'h2D;
		16'hA787: out_word = 8'h44;
		16'hA788: out_word = 8'h4F;
		16'hA789: out_word = 8'hD3;
		16'hA78A: out_word = 8'h20;
		16'hA78B: out_word = 8'h20;
		16'hA78C: out_word = 8'h20;
		16'hA78D: out_word = 8'h20;
		16'hA78E: out_word = 8'h20;
		16'hA78F: out_word = 8'hA0;
		16'hA790: out_word = 8'h05;
		16'hA791: out_word = 8'h00;
		16'hA792: out_word = 8'h42;
		16'hA793: out_word = 8'h27;
		16'hA794: out_word = 8'h01;
		16'hA795: out_word = 8'h51;
		16'hA796: out_word = 8'h28;
		16'hA797: out_word = 8'h02;
		16'hA798: out_word = 8'h11;
		16'hA799: out_word = 8'h28;
		16'hA79A: out_word = 8'h03;
		16'hA79B: out_word = 8'h62;
		16'hA79C: out_word = 8'h28;
		16'hA79D: out_word = 8'h04;
		16'hA79E: out_word = 8'h1C;
		16'hA79F: out_word = 8'h28;
		16'hA7A0: out_word = 8'h06;
		16'hA7A1: out_word = 8'h4F;
		16'hA7A2: out_word = 8'h70;
		16'hA7A3: out_word = 8'h74;
		16'hA7A4: out_word = 8'h69;
		16'hA7A5: out_word = 8'h6F;
		16'hA7A6: out_word = 8'h6E;
		16'hA7A7: out_word = 8'h73;
		16'hA7A8: out_word = 8'h20;
		16'hA7A9: out_word = 8'hFF;
		16'hA7AA: out_word = 8'h31;
		16'hA7AB: out_word = 8'h32;
		16'hA7AC: out_word = 8'h38;
		16'hA7AD: out_word = 8'h20;
		16'hA7AE: out_word = 8'h42;
		16'hA7AF: out_word = 8'h41;
		16'hA7B0: out_word = 8'h53;
		16'hA7B1: out_word = 8'h49;
		16'hA7B2: out_word = 8'hC3;
		16'hA7B3: out_word = 8'h52;
		16'hA7B4: out_word = 8'h65;
		16'hA7B5: out_word = 8'h6E;
		16'hA7B6: out_word = 8'h75;
		16'hA7B7: out_word = 8'h6D;
		16'hA7B8: out_word = 8'h62;
		16'hA7B9: out_word = 8'h65;
		16'hA7BA: out_word = 8'hF2;
		16'hA7BB: out_word = 8'h53;
		16'hA7BC: out_word = 8'h63;
		16'hA7BD: out_word = 8'h72;
		16'hA7BE: out_word = 8'h65;
		16'hA7BF: out_word = 8'h65;
		16'hA7C0: out_word = 8'hEE;
		16'hA7C1: out_word = 8'h50;
		16'hA7C2: out_word = 8'h72;
		16'hA7C3: out_word = 8'h69;
		16'hA7C4: out_word = 8'h6E;
		16'hA7C5: out_word = 8'hF4;
		16'hA7C6: out_word = 8'h45;
		16'hA7C7: out_word = 8'h78;
		16'hA7C8: out_word = 8'h69;
		16'hA7C9: out_word = 8'hF4;
		16'hA7CA: out_word = 8'hA0;
		16'hA7CB: out_word = 8'h02;
		16'hA7CC: out_word = 8'h00;
		16'hA7CD: out_word = 8'h42;
		16'hA7CE: out_word = 8'h27;
		16'hA7CF: out_word = 8'h01;
		16'hA7D0: out_word = 8'h1C;
		16'hA7D1: out_word = 8'h28;
		16'hA7D2: out_word = 8'h03;
		16'hA7D3: out_word = 8'h4F;
		16'hA7D4: out_word = 8'h70;
		16'hA7D5: out_word = 8'h74;
		16'hA7D6: out_word = 8'h69;
		16'hA7D7: out_word = 8'h6F;
		16'hA7D8: out_word = 8'h6E;
		16'hA7D9: out_word = 8'h73;
		16'hA7DA: out_word = 8'h20;
		16'hA7DB: out_word = 8'hFF;
		16'hA7DC: out_word = 8'h43;
		16'hA7DD: out_word = 8'h61;
		16'hA7DE: out_word = 8'h6C;
		16'hA7DF: out_word = 8'h63;
		16'hA7E0: out_word = 8'h75;
		16'hA7E1: out_word = 8'h6C;
		16'hA7E2: out_word = 8'h61;
		16'hA7E3: out_word = 8'h74;
		16'hA7E4: out_word = 8'h6F;
		16'hA7E5: out_word = 8'hF2;
		16'hA7E6: out_word = 8'h45;
		16'hA7E7: out_word = 8'h78;
		16'hA7E8: out_word = 8'h69;
		16'hA7E9: out_word = 8'hF4;
		16'hA7EA: out_word = 8'hA0;
		16'hA7EB: out_word = 8'h16;
		16'hA7EC: out_word = 8'h01;
		16'hA7ED: out_word = 8'h00;
		16'hA7EE: out_word = 8'h10;
		16'hA7EF: out_word = 8'h00;
		16'hA7F0: out_word = 8'h11;
		16'hA7F1: out_word = 8'h07;
		16'hA7F2: out_word = 8'h13;
		16'hA7F3: out_word = 8'h00;
		16'hA7F4: out_word = 8'h54;
		16'hA7F5: out_word = 8'h6F;
		16'hA7F6: out_word = 8'h20;
		16'hA7F7: out_word = 8'h63;
		16'hA7F8: out_word = 8'h61;
		16'hA7F9: out_word = 8'h6E;
		16'hA7FA: out_word = 8'h63;
		16'hA7FB: out_word = 8'h65;
		16'hA7FC: out_word = 8'h6C;
		16'hA7FD: out_word = 8'h20;
		16'hA7FE: out_word = 8'h2D;
		16'hA7FF: out_word = 8'h20;
		16'hA800: out_word = 8'h70;
		16'hA801: out_word = 8'h72;
		16'hA802: out_word = 8'h65;
		16'hA803: out_word = 8'h73;
		16'hA804: out_word = 8'h73;
		16'hA805: out_word = 8'h20;
		16'hA806: out_word = 8'h42;
		16'hA807: out_word = 8'h52;
		16'hA808: out_word = 8'h45;
		16'hA809: out_word = 8'h41;
		16'hA80A: out_word = 8'h4B;
		16'hA80B: out_word = 8'h20;
		16'hA80C: out_word = 8'h74;
		16'hA80D: out_word = 8'h77;
		16'hA80E: out_word = 8'h69;
		16'hA80F: out_word = 8'h63;
		16'hA810: out_word = 8'hE5;
		16'hA811: out_word = 8'hCD;
		16'hA812: out_word = 8'h9B;
		16'hA813: out_word = 8'h26;
		16'hA814: out_word = 8'h18;
		16'hA815: out_word = 8'h5E;
		16'hA816: out_word = 8'hCD;
		16'hA817: out_word = 8'h81;
		16'hA818: out_word = 8'h38;
		16'hA819: out_word = 8'hC3;
		16'hA81A: out_word = 8'hEC;
		16'hA81B: out_word = 8'h3B;
		16'hA81C: out_word = 8'h21;
		16'hA81D: out_word = 8'h0D;
		16'hA81E: out_word = 8'hEC;
		16'hA81F: out_word = 8'hCB;
		16'hA820: out_word = 8'hB6;
		16'hA821: out_word = 8'hCD;
		16'hA822: out_word = 8'hBE;
		16'hA823: out_word = 8'h28;
		16'hA824: out_word = 8'h06;
		16'hA825: out_word = 8'h00;
		16'hA826: out_word = 8'h16;
		16'hA827: out_word = 8'h17;
		16'hA828: out_word = 8'hCD;
		16'hA829: out_word = 8'h5E;
		16'hA82A: out_word = 8'h3B;
		16'hA82B: out_word = 8'hCD;
		16'hA82C: out_word = 8'h20;
		16'hA82D: out_word = 8'h1F;
		16'hA82E: out_word = 8'hC3;
		16'hA82F: out_word = 8'h9F;
		16'hA830: out_word = 8'h25;
		16'hA831: out_word = 8'hCD;
		16'hA832: out_word = 8'h52;
		16'hA833: out_word = 8'h38;
		16'hA834: out_word = 8'h21;
		16'hA835: out_word = 8'h3C;
		16'hA836: out_word = 8'h5C;
		16'hA837: out_word = 8'hCB;
		16'hA838: out_word = 8'hC6;
		16'hA839: out_word = 8'h11;
		16'hA83A: out_word = 8'hEB;
		16'hA83B: out_word = 8'h27;
		16'hA83C: out_word = 8'hCD;
		16'hA83D: out_word = 8'h7D;
		16'hA83E: out_word = 8'h05;
		16'hA83F: out_word = 8'hCB;
		16'hA840: out_word = 8'h86;
		16'hA841: out_word = 8'hCB;
		16'hA842: out_word = 8'hF6;
		16'hA843: out_word = 8'h3E;
		16'hA844: out_word = 8'h07;
		16'hA845: out_word = 8'h32;
		16'hA846: out_word = 8'h0E;
		16'hA847: out_word = 8'hEC;
		16'hA848: out_word = 8'h01;
		16'hA849: out_word = 8'h00;
		16'hA84A: out_word = 8'h00;
		16'hA84B: out_word = 8'hCD;
		16'hA84C: out_word = 8'h2B;
		16'hA84D: out_word = 8'h37;
		16'hA84E: out_word = 8'hC3;
		16'hA84F: out_word = 8'hF1;
		16'hA850: out_word = 8'h1A;
		16'hA851: out_word = 8'hCD;
		16'hA852: out_word = 8'h88;
		16'hA853: out_word = 8'h38;
		16'hA854: out_word = 8'hD4;
		16'hA855: out_word = 8'hE7;
		16'hA856: out_word = 8'h26;
		16'hA857: out_word = 8'h21;
		16'hA858: out_word = 8'h00;
		16'hA859: out_word = 8'h00;
		16'hA85A: out_word = 8'h22;
		16'hA85B: out_word = 8'h49;
		16'hA85C: out_word = 8'h5C;
		16'hA85D: out_word = 8'h22;
		16'hA85E: out_word = 8'h08;
		16'hA85F: out_word = 8'hEC;
		16'hA860: out_word = 8'h18;
		16'hA861: out_word = 8'h03;
		16'hA862: out_word = 8'hCD;
		16'hA863: out_word = 8'h14;
		16'hA864: out_word = 8'h1B;
		16'hA865: out_word = 8'h21;
		16'hA866: out_word = 8'h0D;
		16'hA867: out_word = 8'hEC;
		16'hA868: out_word = 8'hCB;
		16'hA869: out_word = 8'h76;
		16'hA86A: out_word = 8'h20;
		16'hA86B: out_word = 8'h08;
		16'hA86C: out_word = 8'h21;
		16'hA86D: out_word = 8'h3C;
		16'hA86E: out_word = 8'h5C;
		16'hA86F: out_word = 8'hCB;
		16'hA870: out_word = 8'h86;
		16'hA871: out_word = 8'hCD;
		16'hA872: out_word = 8'h48;
		16'hA873: out_word = 8'h38;
		16'hA874: out_word = 8'h21;
		16'hA875: out_word = 8'h0D;
		16'hA876: out_word = 8'hEC;
		16'hA877: out_word = 8'hCB;
		16'hA878: out_word = 8'hAE;
		16'hA879: out_word = 8'hCB;
		16'hA87A: out_word = 8'hA6;
		16'hA87B: out_word = 8'h3E;
		16'hA87C: out_word = 8'h00;
		16'hA87D: out_word = 8'h21;
		16'hA87E: out_word = 8'h90;
		16'hA87F: out_word = 8'h27;
		16'hA880: out_word = 8'h11;
		16'hA881: out_word = 8'hA0;
		16'hA882: out_word = 8'h27;
		16'hA883: out_word = 8'h18;
		16'hA884: out_word = 8'h2C;
		16'hA885: out_word = 8'h21;
		16'hA886: out_word = 8'h0D;
		16'hA887: out_word = 8'hEC;
		16'hA888: out_word = 8'hCB;
		16'hA889: out_word = 8'hEE;
		16'hA88A: out_word = 8'hCB;
		16'hA88B: out_word = 8'hE6;
		16'hA88C: out_word = 8'hCB;
		16'hA88D: out_word = 8'hB6;
		16'hA88E: out_word = 8'hCD;
		16'hA88F: out_word = 8'hBE;
		16'hA890: out_word = 8'h28;
		16'hA891: out_word = 8'hCD;
		16'hA892: out_word = 8'h4D;
		16'hA893: out_word = 8'h38;
		16'hA894: out_word = 8'h3E;
		16'hA895: out_word = 8'h04;
		16'hA896: out_word = 8'h32;
		16'hA897: out_word = 8'h0E;
		16'hA898: out_word = 8'hEC;
		16'hA899: out_word = 8'h21;
		16'hA89A: out_word = 8'h00;
		16'hA89B: out_word = 8'h00;
		16'hA89C: out_word = 8'h22;
		16'hA89D: out_word = 8'h49;
		16'hA89E: out_word = 8'h5C;
		16'hA89F: out_word = 8'hCD;
		16'hA8A0: out_word = 8'h2F;
		16'hA8A1: out_word = 8'h15;
		16'hA8A2: out_word = 8'h01;
		16'hA8A3: out_word = 8'h00;
		16'hA8A4: out_word = 8'h00;
		16'hA8A5: out_word = 8'h78;
		16'hA8A6: out_word = 8'hCD;
		16'hA8A7: out_word = 8'hF8;
		16'hA8A8: out_word = 8'h29;
		16'hA8A9: out_word = 8'h3E;
		16'hA8AA: out_word = 8'h04;
		16'hA8AB: out_word = 8'h21;
		16'hA8AC: out_word = 8'hCB;
		16'hA8AD: out_word = 8'h27;
		16'hA8AE: out_word = 8'h11;
		16'hA8AF: out_word = 8'hD2;
		16'hA8B0: out_word = 8'h27;
		16'hA8B1: out_word = 8'h32;
		16'hA8B2: out_word = 8'h0E;
		16'hA8B3: out_word = 8'hEC;
		16'hA8B4: out_word = 8'h22;
		16'hA8B5: out_word = 8'hEA;
		16'hA8B6: out_word = 8'hF6;
		16'hA8B7: out_word = 8'hED;
		16'hA8B8: out_word = 8'h53;
		16'hA8B9: out_word = 8'hEC;
		16'hA8BA: out_word = 8'hF6;
		16'hA8BB: out_word = 8'hC3;
		16'hA8BC: out_word = 8'h04;
		16'hA8BD: out_word = 8'h26;
		16'hA8BE: out_word = 8'hCD;
		16'hA8BF: out_word = 8'h1F;
		16'hA8C0: out_word = 8'h2E;
		16'hA8C1: out_word = 8'hCD;
		16'hA8C2: out_word = 8'h7F;
		16'hA8C3: out_word = 8'h3A;
		16'hA8C4: out_word = 8'hC3;
		16'hA8C5: out_word = 8'hE8;
		16'hA8C6: out_word = 8'h28;
		16'hA8C7: out_word = 8'h06;
		16'hA8C8: out_word = 8'h00;
		16'hA8C9: out_word = 8'h16;
		16'hA8CA: out_word = 8'h17;
		16'hA8CB: out_word = 8'hCD;
		16'hA8CC: out_word = 8'h5E;
		16'hA8CD: out_word = 8'h3B;
		16'hA8CE: out_word = 8'hC3;
		16'hA8CF: out_word = 8'hAD;
		16'hA8D0: out_word = 8'h25;
		16'hA8D1: out_word = 8'h06;
		16'hA8D2: out_word = 8'h00;
		16'hA8D3: out_word = 8'h00;
		16'hA8D4: out_word = 8'h00;
		16'hA8D5: out_word = 8'h04;
		16'hA8D6: out_word = 8'h10;
		16'hA8D7: out_word = 8'h14;
		16'hA8D8: out_word = 8'h06;
		16'hA8D9: out_word = 8'h00;
		16'hA8DA: out_word = 8'h00;
		16'hA8DB: out_word = 8'h00;
		16'hA8DC: out_word = 8'h00;
		16'hA8DD: out_word = 8'h01;
		16'hA8DE: out_word = 8'h01;
		16'hA8DF: out_word = 8'h21;
		16'hA8E0: out_word = 8'hD8;
		16'hA8E1: out_word = 8'h28;
		16'hA8E2: out_word = 8'h11;
		16'hA8E3: out_word = 8'hEE;
		16'hA8E4: out_word = 8'hF6;
		16'hA8E5: out_word = 8'hC3;
		16'hA8E6: out_word = 8'hBA;
		16'hA8E7: out_word = 8'h3F;
		16'hA8E8: out_word = 8'h21;
		16'hA8E9: out_word = 8'hD1;
		16'hA8EA: out_word = 8'h28;
		16'hA8EB: out_word = 8'h11;
		16'hA8EC: out_word = 8'hEE;
		16'hA8ED: out_word = 8'hF6;
		16'hA8EE: out_word = 8'hC3;
		16'hA8EF: out_word = 8'hBA;
		16'hA8F0: out_word = 8'h3F;
		16'hA8F1: out_word = 8'h21;
		16'hA8F2: out_word = 8'h0D;
		16'hA8F3: out_word = 8'hEC;
		16'hA8F4: out_word = 8'hB7;
		16'hA8F5: out_word = 8'hB7;
		16'hA8F6: out_word = 8'hCB;
		16'hA8F7: out_word = 8'h46;
		16'hA8F8: out_word = 8'hC2;
		16'hA8F9: out_word = 8'hF2;
		16'hA8FA: out_word = 8'h29;
		16'hA8FB: out_word = 8'hCB;
		16'hA8FC: out_word = 8'hBE;
		16'hA8FD: out_word = 8'hCB;
		16'hA8FE: out_word = 8'hDE;
		16'hA8FF: out_word = 8'hE5;
		16'hA900: out_word = 8'hF5;
		16'hA901: out_word = 8'hCD;
		16'hA902: out_word = 8'hEC;
		16'hA903: out_word = 8'h29;
		16'hA904: out_word = 8'hF1;
		16'hA905: out_word = 8'hF5;
		16'hA906: out_word = 8'hCD;
		16'hA907: out_word = 8'h81;
		16'hA908: out_word = 8'h2E;
		16'hA909: out_word = 8'hF1;
		16'hA90A: out_word = 8'h78;
		16'hA90B: out_word = 8'hCD;
		16'hA90C: out_word = 8'h78;
		16'hA90D: out_word = 8'h2B;
		16'hA90E: out_word = 8'hE1;
		16'hA90F: out_word = 8'hCB;
		16'hA910: out_word = 8'hFE;
		16'hA911: out_word = 8'hD2;
		16'hA912: out_word = 8'hF2;
		16'hA913: out_word = 8'h29;
		16'hA914: out_word = 8'h78;
		16'hA915: out_word = 8'hDA;
		16'hA916: out_word = 8'hF8;
		16'hA917: out_word = 8'h29;
		16'hA918: out_word = 8'hC3;
		16'hA919: out_word = 8'hF2;
		16'hA91A: out_word = 8'h29;
		16'hA91B: out_word = 8'h21;
		16'hA91C: out_word = 8'h0D;
		16'hA91D: out_word = 8'hEC;
		16'hA91E: out_word = 8'hCB;
		16'hA91F: out_word = 8'hDE;
		16'hA920: out_word = 8'hCD;
		16'hA921: out_word = 8'hEC;
		16'hA922: out_word = 8'h29;
		16'hA923: out_word = 8'hCD;
		16'hA924: out_word = 8'h12;
		16'hA925: out_word = 8'h2F;
		16'hA926: out_word = 8'h37;
		16'hA927: out_word = 8'h78;
		16'hA928: out_word = 8'hC3;
		16'hA929: out_word = 8'hF8;
		16'hA92A: out_word = 8'h29;
		16'hA92B: out_word = 8'h21;
		16'hA92C: out_word = 8'h0D;
		16'hA92D: out_word = 8'hEC;
		16'hA92E: out_word = 8'hCB;
		16'hA92F: out_word = 8'h86;
		16'hA930: out_word = 8'hCB;
		16'hA931: out_word = 8'hDE;
		16'hA932: out_word = 8'hCD;
		16'hA933: out_word = 8'hEC;
		16'hA934: out_word = 8'h29;
		16'hA935: out_word = 8'hCD;
		16'hA936: out_word = 8'h5B;
		16'hA937: out_word = 8'h2B;
		16'hA938: out_word = 8'h3F;
		16'hA939: out_word = 8'hDA;
		16'hA93A: out_word = 8'hF2;
		16'hA93B: out_word = 8'h29;
		16'hA93C: out_word = 8'hCD;
		16'hA93D: out_word = 8'h12;
		16'hA93E: out_word = 8'h2F;
		16'hA93F: out_word = 8'h37;
		16'hA940: out_word = 8'h78;
		16'hA941: out_word = 8'hC3;
		16'hA942: out_word = 8'hF8;
		16'hA943: out_word = 8'h29;
		16'hA944: out_word = 8'hCD;
		16'hA945: out_word = 8'hEC;
		16'hA946: out_word = 8'h29;
		16'hA947: out_word = 8'hF5;
		16'hA948: out_word = 8'hCD;
		16'hA949: out_word = 8'hB4;
		16'hA94A: out_word = 8'h30;
		16'hA94B: out_word = 8'hC5;
		16'hA94C: out_word = 8'h06;
		16'hA94D: out_word = 8'h00;
		16'hA94E: out_word = 8'hCD;
		16'hA94F: out_word = 8'h41;
		16'hA950: out_word = 8'h2E;
		16'hA951: out_word = 8'hC1;
		16'hA952: out_word = 8'h38;
		16'hA953: out_word = 8'h0A;
		16'hA954: out_word = 8'h21;
		16'hA955: out_word = 8'h20;
		16'hA956: out_word = 8'h00;
		16'hA957: out_word = 8'h19;
		16'hA958: out_word = 8'h7E;
		16'hA959: out_word = 8'h2F;
		16'hA95A: out_word = 8'hE6;
		16'hA95B: out_word = 8'h09;
		16'hA95C: out_word = 8'h28;
		16'hA95D: out_word = 8'h1C;
		16'hA95E: out_word = 8'h3A;
		16'hA95F: out_word = 8'h0D;
		16'hA960: out_word = 8'hEC;
		16'hA961: out_word = 8'hCB;
		16'hA962: out_word = 8'h5F;
		16'hA963: out_word = 8'h28;
		16'hA964: out_word = 8'h05;
		16'hA965: out_word = 8'hCD;
		16'hA966: out_word = 8'h8E;
		16'hA967: out_word = 8'h2C;
		16'hA968: out_word = 8'h30;
		16'hA969: out_word = 8'h15;
		16'hA96A: out_word = 8'hCD;
		16'hA96B: out_word = 8'h4C;
		16'hA96C: out_word = 8'h2C;
		16'hA96D: out_word = 8'hCD;
		16'hA96E: out_word = 8'h78;
		16'hA96F: out_word = 8'h2B;
		16'hA970: out_word = 8'hCD;
		16'hA971: out_word = 8'hCE;
		16'hA972: out_word = 8'h2E;
		16'hA973: out_word = 8'h06;
		16'hA974: out_word = 8'h00;
		16'hA975: out_word = 8'hF1;
		16'hA976: out_word = 8'h37;
		16'hA977: out_word = 8'hC3;
		16'hA978: out_word = 8'hF8;
		16'hA979: out_word = 8'h29;
		16'hA97A: out_word = 8'hF1;
		16'hA97B: out_word = 8'h37;
		16'hA97C: out_word = 8'hC3;
		16'hA97D: out_word = 8'hF2;
		16'hA97E: out_word = 8'h29;
		16'hA97F: out_word = 8'hF1;
		16'hA980: out_word = 8'hC3;
		16'hA981: out_word = 8'hF2;
		16'hA982: out_word = 8'h29;
		16'hA983: out_word = 8'h3A;
		16'hA984: out_word = 8'h0E;
		16'hA985: out_word = 8'hEC;
		16'hA986: out_word = 8'hFE;
		16'hA987: out_word = 8'h04;
		16'hA988: out_word = 8'hC8;
		16'hA989: out_word = 8'hCD;
		16'hA98A: out_word = 8'hEC;
		16'hA98B: out_word = 8'h29;
		16'hA98C: out_word = 8'h21;
		16'hA98D: out_word = 8'h00;
		16'hA98E: out_word = 8'h00;
		16'hA98F: out_word = 8'hCD;
		16'hA990: out_word = 8'h20;
		16'hA991: out_word = 8'h1F;
		16'hA992: out_word = 8'hEF;
		16'hA993: out_word = 8'h6E;
		16'hA994: out_word = 8'h19;
		16'hA995: out_word = 8'hEF;
		16'hA996: out_word = 8'h95;
		16'hA997: out_word = 8'h16;
		16'hA998: out_word = 8'hCD;
		16'hA999: out_word = 8'h45;
		16'hA99A: out_word = 8'h1F;
		16'hA99B: out_word = 8'hED;
		16'hA99C: out_word = 8'h53;
		16'hA99D: out_word = 8'h49;
		16'hA99E: out_word = 8'h5C;
		16'hA99F: out_word = 8'h3E;
		16'hA9A0: out_word = 8'h0F;
		16'hA9A1: out_word = 8'hCD;
		16'hA9A2: out_word = 8'h96;
		16'hA9A3: out_word = 8'h3A;
		16'hA9A4: out_word = 8'hCD;
		16'hA9A5: out_word = 8'h2F;
		16'hA9A6: out_word = 8'h15;
		16'hA9A7: out_word = 8'h37;
		16'hA9A8: out_word = 8'hC3;
		16'hA9A9: out_word = 8'hF2;
		16'hA9AA: out_word = 8'h29;
		16'hA9AB: out_word = 8'h3A;
		16'hA9AC: out_word = 8'h0E;
		16'hA9AD: out_word = 8'hEC;
		16'hA9AE: out_word = 8'hFE;
		16'hA9AF: out_word = 8'h04;
		16'hA9B0: out_word = 8'hC8;
		16'hA9B1: out_word = 8'hCD;
		16'hA9B2: out_word = 8'hEC;
		16'hA9B3: out_word = 8'h29;
		16'hA9B4: out_word = 8'h21;
		16'hA9B5: out_word = 8'h0F;
		16'hA9B6: out_word = 8'h27;
		16'hA9B7: out_word = 8'hCD;
		16'hA9B8: out_word = 8'h20;
		16'hA9B9: out_word = 8'h1F;
		16'hA9BA: out_word = 8'hEF;
		16'hA9BB: out_word = 8'h6E;
		16'hA9BC: out_word = 8'h19;
		16'hA9BD: out_word = 8'hEB;
		16'hA9BE: out_word = 8'hEF;
		16'hA9BF: out_word = 8'h95;
		16'hA9C0: out_word = 8'h16;
		16'hA9C1: out_word = 8'hCD;
		16'hA9C2: out_word = 8'h45;
		16'hA9C3: out_word = 8'h1F;
		16'hA9C4: out_word = 8'hED;
		16'hA9C5: out_word = 8'h53;
		16'hA9C6: out_word = 8'h49;
		16'hA9C7: out_word = 8'h5C;
		16'hA9C8: out_word = 8'h3E;
		16'hA9C9: out_word = 8'h0F;
		16'hA9CA: out_word = 8'hCD;
		16'hA9CB: out_word = 8'h96;
		16'hA9CC: out_word = 8'h3A;
		16'hA9CD: out_word = 8'hCD;
		16'hA9CE: out_word = 8'h2F;
		16'hA9CF: out_word = 8'h15;
		16'hA9D0: out_word = 8'h37;
		16'hA9D1: out_word = 8'hC3;
		16'hA9D2: out_word = 8'hF2;
		16'hA9D3: out_word = 8'h29;
		16'hA9D4: out_word = 8'hCD;
		16'hA9D5: out_word = 8'hEC;
		16'hA9D6: out_word = 8'h29;
		16'hA9D7: out_word = 8'hCD;
		16'hA9D8: out_word = 8'hEA;
		16'hA9D9: out_word = 8'h2B;
		16'hA9DA: out_word = 8'hD2;
		16'hA9DB: out_word = 8'hF2;
		16'hA9DC: out_word = 8'h29;
		16'hA9DD: out_word = 8'h78;
		16'hA9DE: out_word = 8'hC3;
		16'hA9DF: out_word = 8'hF8;
		16'hA9E0: out_word = 8'h29;
		16'hA9E1: out_word = 8'hCD;
		16'hA9E2: out_word = 8'hEC;
		16'hA9E3: out_word = 8'h29;
		16'hA9E4: out_word = 8'hCD;
		16'hA9E5: out_word = 8'h09;
		16'hA9E6: out_word = 8'h2C;
		16'hA9E7: out_word = 8'h30;
		16'hA9E8: out_word = 8'h09;
		16'hA9E9: out_word = 8'h78;
		16'hA9EA: out_word = 8'h18;
		16'hA9EB: out_word = 8'h0C;
		16'hA9EC: out_word = 8'hCD;
		16'hA9ED: out_word = 8'h07;
		16'hA9EE: out_word = 8'h2A;
		16'hA9EF: out_word = 8'hC3;
		16'hA9F0: out_word = 8'h4F;
		16'hA9F1: out_word = 8'h36;
		16'hA9F2: out_word = 8'hCD;
		16'hA9F3: out_word = 8'h07;
		16'hA9F4: out_word = 8'h2A;
		16'hA9F5: out_word = 8'hC3;
		16'hA9F6: out_word = 8'h40;
		16'hA9F7: out_word = 8'h36;
		16'hA9F8: out_word = 8'hCD;
		16'hA9F9: out_word = 8'h11;
		16'hA9FA: out_word = 8'h2A;
		16'hA9FB: out_word = 8'hF5;
		16'hA9FC: out_word = 8'hC5;
		16'hA9FD: out_word = 8'h3E;
		16'hA9FE: out_word = 8'h0F;
		16'hA9FF: out_word = 8'hCD;
		16'hAA00: out_word = 8'h96;
		16'hAA01: out_word = 8'h3A;
		16'hAA02: out_word = 8'hC1;
		16'hAA03: out_word = 8'hF1;
		16'hAA04: out_word = 8'hC3;
		16'hAA05: out_word = 8'h40;
		16'hAA06: out_word = 8'h36;
		16'hAA07: out_word = 8'h21;
		16'hAA08: out_word = 8'hEE;
		16'hAA09: out_word = 8'hF6;
		16'hAA0A: out_word = 8'h4E;
		16'hAA0B: out_word = 8'h23;
		16'hAA0C: out_word = 8'h46;
		16'hAA0D: out_word = 8'h23;
		16'hAA0E: out_word = 8'h7E;
		16'hAA0F: out_word = 8'h23;
		16'hAA10: out_word = 8'hC9;
		16'hAA11: out_word = 8'h21;
		16'hAA12: out_word = 8'hEE;
		16'hAA13: out_word = 8'hF6;
		16'hAA14: out_word = 8'h71;
		16'hAA15: out_word = 8'h23;
		16'hAA16: out_word = 8'h70;
		16'hAA17: out_word = 8'h23;
		16'hAA18: out_word = 8'h77;
		16'hAA19: out_word = 8'hC9;
		16'hAA1A: out_word = 8'hE5;
		16'hAA1B: out_word = 8'hCD;
		16'hAA1C: out_word = 8'hB4;
		16'hAA1D: out_word = 8'h30;
		16'hAA1E: out_word = 8'h26;
		16'hAA1F: out_word = 8'h00;
		16'hAA20: out_word = 8'h68;
		16'hAA21: out_word = 8'h19;
		16'hAA22: out_word = 8'h7E;
		16'hAA23: out_word = 8'hE1;
		16'hAA24: out_word = 8'hC9;
		16'hAA25: out_word = 8'hCD;
		16'hAA26: out_word = 8'hEC;
		16'hAA27: out_word = 8'h29;
		16'hAA28: out_word = 8'h5F;
		16'hAA29: out_word = 8'h16;
		16'hAA2A: out_word = 8'h0A;
		16'hAA2B: out_word = 8'hD5;
		16'hAA2C: out_word = 8'hCD;
		16'hAA2D: out_word = 8'h30;
		16'hAA2E: out_word = 8'h2B;
		16'hAA2F: out_word = 8'hD1;
		16'hAA30: out_word = 8'h30;
		16'hAA31: out_word = 8'hC0;
		16'hAA32: out_word = 8'h7B;
		16'hAA33: out_word = 8'hCD;
		16'hAA34: out_word = 8'h11;
		16'hAA35: out_word = 8'h2A;
		16'hAA36: out_word = 8'h43;
		16'hAA37: out_word = 8'hCD;
		16'hAA38: out_word = 8'hF9;
		16'hAA39: out_word = 8'h2A;
		16'hAA3A: out_word = 8'h30;
		16'hAA3B: out_word = 8'h06;
		16'hAA3C: out_word = 8'h15;
		16'hAA3D: out_word = 8'h20;
		16'hAA3E: out_word = 8'hEC;
		16'hAA3F: out_word = 8'h7B;
		16'hAA40: out_word = 8'h38;
		16'hAA41: out_word = 8'hB6;
		16'hAA42: out_word = 8'hD5;
		16'hAA43: out_word = 8'hCD;
		16'hAA44: out_word = 8'h0B;
		16'hAA45: out_word = 8'h2B;
		16'hAA46: out_word = 8'hD1;
		16'hAA47: out_word = 8'h43;
		16'hAA48: out_word = 8'hCD;
		16'hAA49: out_word = 8'hF9;
		16'hAA4A: out_word = 8'h2A;
		16'hAA4B: out_word = 8'h7B;
		16'hAA4C: out_word = 8'hB7;
		16'hAA4D: out_word = 8'h18;
		16'hAA4E: out_word = 8'hA9;
		16'hAA4F: out_word = 8'hCD;
		16'hAA50: out_word = 8'hEC;
		16'hAA51: out_word = 8'h29;
		16'hAA52: out_word = 8'h5F;
		16'hAA53: out_word = 8'h16;
		16'hAA54: out_word = 8'h0A;
		16'hAA55: out_word = 8'hD5;
		16'hAA56: out_word = 8'hCD;
		16'hAA57: out_word = 8'h0B;
		16'hAA58: out_word = 8'h2B;
		16'hAA59: out_word = 8'hD1;
		16'hAA5A: out_word = 8'h30;
		16'hAA5B: out_word = 8'h96;
		16'hAA5C: out_word = 8'h7B;
		16'hAA5D: out_word = 8'hCD;
		16'hAA5E: out_word = 8'h11;
		16'hAA5F: out_word = 8'h2A;
		16'hAA60: out_word = 8'h43;
		16'hAA61: out_word = 8'hCD;
		16'hAA62: out_word = 8'h02;
		16'hAA63: out_word = 8'h2B;
		16'hAA64: out_word = 8'h30;
		16'hAA65: out_word = 8'h07;
		16'hAA66: out_word = 8'h15;
		16'hAA67: out_word = 8'h20;
		16'hAA68: out_word = 8'hEC;
		16'hAA69: out_word = 8'h7B;
		16'hAA6A: out_word = 8'hDA;
		16'hAA6B: out_word = 8'hF8;
		16'hAA6C: out_word = 8'h29;
		16'hAA6D: out_word = 8'hF5;
		16'hAA6E: out_word = 8'hCD;
		16'hAA6F: out_word = 8'h30;
		16'hAA70: out_word = 8'h2B;
		16'hAA71: out_word = 8'h06;
		16'hAA72: out_word = 8'h00;
		16'hAA73: out_word = 8'hCD;
		16'hAA74: out_word = 8'hD4;
		16'hAA75: out_word = 8'h2B;
		16'hAA76: out_word = 8'hF1;
		16'hAA77: out_word = 8'hC3;
		16'hAA78: out_word = 8'hF8;
		16'hAA79: out_word = 8'h29;
		16'hAA7A: out_word = 8'hCD;
		16'hAA7B: out_word = 8'hEC;
		16'hAA7C: out_word = 8'h29;
		16'hAA7D: out_word = 8'hCD;
		16'hAA7E: out_word = 8'h4C;
		16'hAA7F: out_word = 8'h2C;
		16'hAA80: out_word = 8'hD2;
		16'hAA81: out_word = 8'hF2;
		16'hAA82: out_word = 8'h29;
		16'hAA83: out_word = 8'h78;
		16'hAA84: out_word = 8'hC3;
		16'hAA85: out_word = 8'hF8;
		16'hAA86: out_word = 8'h29;
		16'hAA87: out_word = 8'hCD;
		16'hAA88: out_word = 8'hEC;
		16'hAA89: out_word = 8'h29;
		16'hAA8A: out_word = 8'hCD;
		16'hAA8B: out_word = 8'h31;
		16'hAA8C: out_word = 8'h2C;
		16'hAA8D: out_word = 8'hD2;
		16'hAA8E: out_word = 8'hF2;
		16'hAA8F: out_word = 8'h29;
		16'hAA90: out_word = 8'h78;
		16'hAA91: out_word = 8'hC3;
		16'hAA92: out_word = 8'hF8;
		16'hAA93: out_word = 8'h29;
		16'hAA94: out_word = 8'hCD;
		16'hAA95: out_word = 8'hEC;
		16'hAA96: out_word = 8'h29;
		16'hAA97: out_word = 8'h5F;
		16'hAA98: out_word = 8'hD5;
		16'hAA99: out_word = 8'hCD;
		16'hAA9A: out_word = 8'h0B;
		16'hAA9B: out_word = 8'h2B;
		16'hAA9C: out_word = 8'hD1;
		16'hAA9D: out_word = 8'hD2;
		16'hAA9E: out_word = 8'hF2;
		16'hAA9F: out_word = 8'h29;
		16'hAAA0: out_word = 8'h43;
		16'hAAA1: out_word = 8'hCD;
		16'hAAA2: out_word = 8'h02;
		16'hAAA3: out_word = 8'h2B;
		16'hAAA4: out_word = 8'h7B;
		16'hAAA5: out_word = 8'hDA;
		16'hAAA6: out_word = 8'hF8;
		16'hAAA7: out_word = 8'h29;
		16'hAAA8: out_word = 8'hF5;
		16'hAAA9: out_word = 8'hCD;
		16'hAAAA: out_word = 8'h30;
		16'hAAAB: out_word = 8'h2B;
		16'hAAAC: out_word = 8'h06;
		16'hAAAD: out_word = 8'h00;
		16'hAAAE: out_word = 8'hCD;
		16'hAAAF: out_word = 8'hF9;
		16'hAAB0: out_word = 8'h2A;
		16'hAAB1: out_word = 8'hF1;
		16'hAAB2: out_word = 8'hC3;
		16'hAAB3: out_word = 8'hF8;
		16'hAAB4: out_word = 8'h29;
		16'hAAB5: out_word = 8'hCD;
		16'hAAB6: out_word = 8'hEC;
		16'hAAB7: out_word = 8'h29;
		16'hAAB8: out_word = 8'h5F;
		16'hAAB9: out_word = 8'hD5;
		16'hAABA: out_word = 8'hCD;
		16'hAABB: out_word = 8'h30;
		16'hAABC: out_word = 8'h2B;
		16'hAABD: out_word = 8'hD1;
		16'hAABE: out_word = 8'hD2;
		16'hAABF: out_word = 8'hF2;
		16'hAAC0: out_word = 8'h29;
		16'hAAC1: out_word = 8'h43;
		16'hAAC2: out_word = 8'hCD;
		16'hAAC3: out_word = 8'h02;
		16'hAAC4: out_word = 8'h2B;
		16'hAAC5: out_word = 8'h7B;
		16'hAAC6: out_word = 8'hDA;
		16'hAAC7: out_word = 8'hF8;
		16'hAAC8: out_word = 8'h29;
		16'hAAC9: out_word = 8'hD5;
		16'hAACA: out_word = 8'hCD;
		16'hAACB: out_word = 8'h0B;
		16'hAACC: out_word = 8'h2B;
		16'hAACD: out_word = 8'hD1;
		16'hAACE: out_word = 8'h43;
		16'hAACF: out_word = 8'hCD;
		16'hAAD0: out_word = 8'hF9;
		16'hAAD1: out_word = 8'h2A;
		16'hAAD2: out_word = 8'h7B;
		16'hAAD3: out_word = 8'hB7;
		16'hAAD4: out_word = 8'hC3;
		16'hAAD5: out_word = 8'hF8;
		16'hAAD6: out_word = 8'h29;
		16'hAAD7: out_word = 8'hCD;
		16'hAAD8: out_word = 8'hEC;
		16'hAAD9: out_word = 8'h29;
		16'hAADA: out_word = 8'hCD;
		16'hAADB: out_word = 8'h5B;
		16'hAADC: out_word = 8'h2B;
		16'hAADD: out_word = 8'hDA;
		16'hAADE: out_word = 8'hF8;
		16'hAADF: out_word = 8'h29;
		16'hAAE0: out_word = 8'hC3;
		16'hAAE1: out_word = 8'hF2;
		16'hAAE2: out_word = 8'h29;
		16'hAAE3: out_word = 8'hCD;
		16'hAAE4: out_word = 8'hEC;
		16'hAAE5: out_word = 8'h29;
		16'hAAE6: out_word = 8'hCD;
		16'hAAE7: out_word = 8'h78;
		16'hAAE8: out_word = 8'h2B;
		16'hAAE9: out_word = 8'hDA;
		16'hAAEA: out_word = 8'hF8;
		16'hAAEB: out_word = 8'h29;
		16'hAAEC: out_word = 8'hF5;
		16'hAAED: out_word = 8'hCD;
		16'hAAEE: out_word = 8'h0B;
		16'hAAEF: out_word = 8'h2B;
		16'hAAF0: out_word = 8'h06;
		16'hAAF1: out_word = 8'h1F;
		16'hAAF2: out_word = 8'hCD;
		16'hAAF3: out_word = 8'hDF;
		16'hAAF4: out_word = 8'h2B;
		16'hAAF5: out_word = 8'hF1;
		16'hAAF6: out_word = 8'hC3;
		16'hAAF7: out_word = 8'hF8;
		16'hAAF8: out_word = 8'h29;
		16'hAAF9: out_word = 8'hD5;
		16'hAAFA: out_word = 8'hCD;
		16'hAAFB: out_word = 8'hD4;
		16'hAAFC: out_word = 8'h2B;
		16'hAAFD: out_word = 8'hD4;
		16'hAAFE: out_word = 8'hDF;
		16'hAAFF: out_word = 8'h2B;
		16'hAB00: out_word = 8'hD1;
		16'hAB01: out_word = 8'hC9;
		16'hAB02: out_word = 8'hD5;
		16'hAB03: out_word = 8'hCD;
		16'hAB04: out_word = 8'hDF;
		16'hAB05: out_word = 8'h2B;
		16'hAB06: out_word = 8'hD4;
		16'hAB07: out_word = 8'hD4;
		16'hAB08: out_word = 8'h2B;
		16'hAB09: out_word = 8'hD1;
		16'hAB0A: out_word = 8'hC9;
		16'hAB0B: out_word = 8'hCD;
		16'hAB0C: out_word = 8'h7C;
		16'hAB0D: out_word = 8'h2C;
		16'hAB0E: out_word = 8'h30;
		16'hAB0F: out_word = 8'h1F;
		16'hAB10: out_word = 8'hC5;
		16'hAB11: out_word = 8'hCD;
		16'hAB12: out_word = 8'hB4;
		16'hAB13: out_word = 8'h30;
		16'hAB14: out_word = 8'h06;
		16'hAB15: out_word = 8'h00;
		16'hAB16: out_word = 8'hCD;
		16'hAB17: out_word = 8'h41;
		16'hAB18: out_word = 8'h2E;
		16'hAB19: out_word = 8'hD4;
		16'hAB1A: out_word = 8'h80;
		16'hAB1B: out_word = 8'h2F;
		16'hAB1C: out_word = 8'hC1;
		16'hAB1D: out_word = 8'h21;
		16'hAB1E: out_word = 8'hF1;
		16'hAB1F: out_word = 8'hF6;
		16'hAB20: out_word = 8'h7E;
		16'hAB21: out_word = 8'hB9;
		16'hAB22: out_word = 8'h38;
		16'hAB23: out_word = 8'h09;
		16'hAB24: out_word = 8'hC5;
		16'hAB25: out_word = 8'hCD;
		16'hAB26: out_word = 8'h6F;
		16'hAB27: out_word = 8'h16;
		16'hAB28: out_word = 8'hC1;
		16'hAB29: out_word = 8'hD8;
		16'hAB2A: out_word = 8'h79;
		16'hAB2B: out_word = 8'hB7;
		16'hAB2C: out_word = 8'hC8;
		16'hAB2D: out_word = 8'h0D;
		16'hAB2E: out_word = 8'h37;
		16'hAB2F: out_word = 8'hC9;
		16'hAB30: out_word = 8'hC5;
		16'hAB31: out_word = 8'hCD;
		16'hAB32: out_word = 8'hB4;
		16'hAB33: out_word = 8'h30;
		16'hAB34: out_word = 8'h06;
		16'hAB35: out_word = 8'h00;
		16'hAB36: out_word = 8'hCD;
		16'hAB37: out_word = 8'h41;
		16'hAB38: out_word = 8'h2E;
		16'hAB39: out_word = 8'hC1;
		16'hAB3A: out_word = 8'h38;
		16'hAB3B: out_word = 8'h03;
		16'hAB3C: out_word = 8'hC3;
		16'hAB3D: out_word = 8'h80;
		16'hAB3E: out_word = 8'h2F;
		16'hAB3F: out_word = 8'hCD;
		16'hAB40: out_word = 8'h68;
		16'hAB41: out_word = 8'h2C;
		16'hAB42: out_word = 8'h30;
		16'hAB43: out_word = 8'h16;
		16'hAB44: out_word = 8'h21;
		16'hAB45: out_word = 8'hF1;
		16'hAB46: out_word = 8'hF6;
		16'hAB47: out_word = 8'h23;
		16'hAB48: out_word = 8'h79;
		16'hAB49: out_word = 8'hBE;
		16'hAB4A: out_word = 8'h38;
		16'hAB4B: out_word = 8'h0C;
		16'hAB4C: out_word = 8'hC5;
		16'hAB4D: out_word = 8'hE5;
		16'hAB4E: out_word = 8'hCD;
		16'hAB4F: out_word = 8'h39;
		16'hAB50: out_word = 8'h16;
		16'hAB51: out_word = 8'hE1;
		16'hAB52: out_word = 8'hC1;
		16'hAB53: out_word = 8'hD8;
		16'hAB54: out_word = 8'h23;
		16'hAB55: out_word = 8'h7E;
		16'hAB56: out_word = 8'hB9;
		16'hAB57: out_word = 8'hC8;
		16'hAB58: out_word = 8'h0C;
		16'hAB59: out_word = 8'h37;
		16'hAB5A: out_word = 8'hC9;
		16'hAB5B: out_word = 8'h57;
		16'hAB5C: out_word = 8'h05;
		16'hAB5D: out_word = 8'hFA;
		16'hAB5E: out_word = 8'h66;
		16'hAB5F: out_word = 8'h2B;
		16'hAB60: out_word = 8'h58;
		16'hAB61: out_word = 8'hCD;
		16'hAB62: out_word = 8'hDF;
		16'hAB63: out_word = 8'h2B;
		16'hAB64: out_word = 8'h7B;
		16'hAB65: out_word = 8'hD8;
		16'hAB66: out_word = 8'hD5;
		16'hAB67: out_word = 8'hCD;
		16'hAB68: out_word = 8'h0B;
		16'hAB69: out_word = 8'h2B;
		16'hAB6A: out_word = 8'hD1;
		16'hAB6B: out_word = 8'h7B;
		16'hAB6C: out_word = 8'hD0;
		16'hAB6D: out_word = 8'h06;
		16'hAB6E: out_word = 8'h1F;
		16'hAB6F: out_word = 8'hCD;
		16'hAB70: out_word = 8'hDF;
		16'hAB71: out_word = 8'h2B;
		16'hAB72: out_word = 8'h78;
		16'hAB73: out_word = 8'hD8;
		16'hAB74: out_word = 8'h7A;
		16'hAB75: out_word = 8'h06;
		16'hAB76: out_word = 8'h00;
		16'hAB77: out_word = 8'hC9;
		16'hAB78: out_word = 8'h57;
		16'hAB79: out_word = 8'h04;
		16'hAB7A: out_word = 8'h3E;
		16'hAB7B: out_word = 8'h1F;
		16'hAB7C: out_word = 8'hB8;
		16'hAB7D: out_word = 8'h38;
		16'hAB7E: out_word = 8'h06;
		16'hAB7F: out_word = 8'h58;
		16'hAB80: out_word = 8'hCD;
		16'hAB81: out_word = 8'hD4;
		16'hAB82: out_word = 8'h2B;
		16'hAB83: out_word = 8'h7B;
		16'hAB84: out_word = 8'hD8;
		16'hAB85: out_word = 8'h05;
		16'hAB86: out_word = 8'hC5;
		16'hAB87: out_word = 8'hE5;
		16'hAB88: out_word = 8'h21;
		16'hAB89: out_word = 8'h0D;
		16'hAB8A: out_word = 8'hEC;
		16'hAB8B: out_word = 8'hCB;
		16'hAB8C: out_word = 8'h7E;
		16'hAB8D: out_word = 8'h20;
		16'hAB8E: out_word = 8'h31;
		16'hAB8F: out_word = 8'hCD;
		16'hAB90: out_word = 8'hB4;
		16'hAB91: out_word = 8'h30;
		16'hAB92: out_word = 8'h21;
		16'hAB93: out_word = 8'h20;
		16'hAB94: out_word = 8'h00;
		16'hAB95: out_word = 8'h19;
		16'hAB96: out_word = 8'h7E;
		16'hAB97: out_word = 8'hCB;
		16'hAB98: out_word = 8'h4F;
		16'hAB99: out_word = 8'h20;
		16'hAB9A: out_word = 8'h25;
		16'hAB9B: out_word = 8'hCB;
		16'hAB9C: out_word = 8'hCE;
		16'hAB9D: out_word = 8'hCB;
		16'hAB9E: out_word = 8'h9E;
		16'hAB9F: out_word = 8'h21;
		16'hABA0: out_word = 8'h23;
		16'hABA1: out_word = 8'h00;
		16'hABA2: out_word = 8'h19;
		16'hABA3: out_word = 8'hEB;
		16'hABA4: out_word = 8'hE1;
		16'hABA5: out_word = 8'hC1;
		16'hABA6: out_word = 8'hF5;
		16'hABA7: out_word = 8'hCD;
		16'hABA8: out_word = 8'h30;
		16'hABA9: out_word = 8'h2B;
		16'hABAA: out_word = 8'hF1;
		16'hABAB: out_word = 8'hCD;
		16'hABAC: out_word = 8'hB4;
		16'hABAD: out_word = 8'h30;
		16'hABAE: out_word = 8'h21;
		16'hABAF: out_word = 8'h23;
		16'hABB0: out_word = 8'h00;
		16'hABB1: out_word = 8'h19;
		16'hABB2: out_word = 8'hEB;
		16'hABB3: out_word = 8'hCB;
		16'hABB4: out_word = 8'h87;
		16'hABB5: out_word = 8'hCB;
		16'hABB6: out_word = 8'hDF;
		16'hABB7: out_word = 8'hCD;
		16'hABB8: out_word = 8'hD3;
		16'hABB9: out_word = 8'h2E;
		16'hABBA: out_word = 8'hCD;
		16'hABBB: out_word = 8'hF4;
		16'hABBC: out_word = 8'h35;
		16'hABBD: out_word = 8'h78;
		16'hABBE: out_word = 8'h37;
		16'hABBF: out_word = 8'hC9;
		16'hABC0: out_word = 8'hE1;
		16'hABC1: out_word = 8'hC1;
		16'hABC2: out_word = 8'hD5;
		16'hABC3: out_word = 8'hCD;
		16'hABC4: out_word = 8'h30;
		16'hABC5: out_word = 8'h2B;
		16'hABC6: out_word = 8'hD1;
		16'hABC7: out_word = 8'h78;
		16'hABC8: out_word = 8'hD0;
		16'hABC9: out_word = 8'h06;
		16'hABCA: out_word = 8'h00;
		16'hABCB: out_word = 8'hCD;
		16'hABCC: out_word = 8'hD4;
		16'hABCD: out_word = 8'h2B;
		16'hABCE: out_word = 8'h78;
		16'hABCF: out_word = 8'hD8;
		16'hABD0: out_word = 8'h7B;
		16'hABD1: out_word = 8'h06;
		16'hABD2: out_word = 8'h00;
		16'hABD3: out_word = 8'hC9;
		16'hABD4: out_word = 8'hD5;
		16'hABD5: out_word = 8'hE5;
		16'hABD6: out_word = 8'hCD;
		16'hABD7: out_word = 8'hB4;
		16'hABD8: out_word = 8'h30;
		16'hABD9: out_word = 8'hCD;
		16'hABDA: out_word = 8'h41;
		16'hABDB: out_word = 8'h2E;
		16'hABDC: out_word = 8'hC3;
		16'hABDD: out_word = 8'h65;
		16'hABDE: out_word = 8'h2C;
		16'hABDF: out_word = 8'hD5;
		16'hABE0: out_word = 8'hE5;
		16'hABE1: out_word = 8'hCD;
		16'hABE2: out_word = 8'hB4;
		16'hABE3: out_word = 8'h30;
		16'hABE4: out_word = 8'hCD;
		16'hABE5: out_word = 8'h63;
		16'hABE6: out_word = 8'h2E;
		16'hABE7: out_word = 8'hC3;
		16'hABE8: out_word = 8'h65;
		16'hABE9: out_word = 8'h2C;
		16'hABEA: out_word = 8'hD5;
		16'hABEB: out_word = 8'hE5;
		16'hABEC: out_word = 8'hCD;
		16'hABED: out_word = 8'h5B;
		16'hABEE: out_word = 8'h2B;
		16'hABEF: out_word = 8'h30;
		16'hABF0: out_word = 8'h16;
		16'hABF1: out_word = 8'hCD;
		16'hABF2: out_word = 8'h1A;
		16'hABF3: out_word = 8'h2A;
		16'hABF4: out_word = 8'hFE;
		16'hABF5: out_word = 8'h20;
		16'hABF6: out_word = 8'h28;
		16'hABF7: out_word = 8'hF4;
		16'hABF8: out_word = 8'hCD;
		16'hABF9: out_word = 8'h5B;
		16'hABFA: out_word = 8'h2B;
		16'hABFB: out_word = 8'h30;
		16'hABFC: out_word = 8'h0A;
		16'hABFD: out_word = 8'hCD;
		16'hABFE: out_word = 8'h1A;
		16'hABFF: out_word = 8'h2A;
		16'hAC00: out_word = 8'hFE;
		16'hAC01: out_word = 8'h20;
		16'hAC02: out_word = 8'h20;
		16'hAC03: out_word = 8'hF4;
		16'hAC04: out_word = 8'hCD;
		16'hAC05: out_word = 8'h78;
		16'hAC06: out_word = 8'h2B;
		16'hAC07: out_word = 8'h18;
		16'hAC08: out_word = 8'h5C;
		16'hAC09: out_word = 8'hD5;
		16'hAC0A: out_word = 8'hE5;
		16'hAC0B: out_word = 8'hCD;
		16'hAC0C: out_word = 8'h78;
		16'hAC0D: out_word = 8'h2B;
		16'hAC0E: out_word = 8'h30;
		16'hAC0F: out_word = 8'h1B;
		16'hAC10: out_word = 8'hCD;
		16'hAC11: out_word = 8'h1A;
		16'hAC12: out_word = 8'h2A;
		16'hAC13: out_word = 8'hFE;
		16'hAC14: out_word = 8'h20;
		16'hAC15: out_word = 8'h20;
		16'hAC16: out_word = 8'hF4;
		16'hAC17: out_word = 8'hCD;
		16'hAC18: out_word = 8'h78;
		16'hAC19: out_word = 8'h2B;
		16'hAC1A: out_word = 8'h30;
		16'hAC1B: out_word = 8'h0F;
		16'hAC1C: out_word = 8'hCD;
		16'hAC1D: out_word = 8'h41;
		16'hAC1E: out_word = 8'h2E;
		16'hAC1F: out_word = 8'h30;
		16'hAC20: out_word = 8'h0A;
		16'hAC21: out_word = 8'hCD;
		16'hAC22: out_word = 8'h1A;
		16'hAC23: out_word = 8'h2A;
		16'hAC24: out_word = 8'hFE;
		16'hAC25: out_word = 8'h20;
		16'hAC26: out_word = 8'h28;
		16'hAC27: out_word = 8'hEF;
		16'hAC28: out_word = 8'h37;
		16'hAC29: out_word = 8'h18;
		16'hAC2A: out_word = 8'h3A;
		16'hAC2B: out_word = 8'hD4;
		16'hAC2C: out_word = 8'h5B;
		16'hAC2D: out_word = 8'h2B;
		16'hAC2E: out_word = 8'hB7;
		16'hAC2F: out_word = 8'h18;
		16'hAC30: out_word = 8'h34;
		16'hAC31: out_word = 8'hD5;
		16'hAC32: out_word = 8'hE5;
		16'hAC33: out_word = 8'hCD;
		16'hAC34: out_word = 8'hB4;
		16'hAC35: out_word = 8'h30;
		16'hAC36: out_word = 8'h21;
		16'hAC37: out_word = 8'h20;
		16'hAC38: out_word = 8'h00;
		16'hAC39: out_word = 8'h19;
		16'hAC3A: out_word = 8'hCB;
		16'hAC3B: out_word = 8'h46;
		16'hAC3C: out_word = 8'h20;
		16'hAC3D: out_word = 8'h07;
		16'hAC3E: out_word = 8'hCD;
		16'hAC3F: out_word = 8'h0B;
		16'hAC40: out_word = 8'h2B;
		16'hAC41: out_word = 8'h38;
		16'hAC42: out_word = 8'hF0;
		16'hAC43: out_word = 8'h18;
		16'hAC44: out_word = 8'h20;
		16'hAC45: out_word = 8'h06;
		16'hAC46: out_word = 8'h00;
		16'hAC47: out_word = 8'hCD;
		16'hAC48: out_word = 8'hD4;
		16'hAC49: out_word = 8'h2B;
		16'hAC4A: out_word = 8'h18;
		16'hAC4B: out_word = 8'h19;
		16'hAC4C: out_word = 8'hD5;
		16'hAC4D: out_word = 8'hE5;
		16'hAC4E: out_word = 8'hCD;
		16'hAC4F: out_word = 8'hB4;
		16'hAC50: out_word = 8'h30;
		16'hAC51: out_word = 8'h21;
		16'hAC52: out_word = 8'h20;
		16'hAC53: out_word = 8'h00;
		16'hAC54: out_word = 8'h19;
		16'hAC55: out_word = 8'hCB;
		16'hAC56: out_word = 8'h5E;
		16'hAC57: out_word = 8'h20;
		16'hAC58: out_word = 8'h07;
		16'hAC59: out_word = 8'hCD;
		16'hAC5A: out_word = 8'h30;
		16'hAC5B: out_word = 8'h2B;
		16'hAC5C: out_word = 8'h38;
		16'hAC5D: out_word = 8'hF0;
		16'hAC5E: out_word = 8'h18;
		16'hAC5F: out_word = 8'h05;
		16'hAC60: out_word = 8'h06;
		16'hAC61: out_word = 8'h1F;
		16'hAC62: out_word = 8'hCD;
		16'hAC63: out_word = 8'hDF;
		16'hAC64: out_word = 8'h2B;
		16'hAC65: out_word = 8'hE1;
		16'hAC66: out_word = 8'hD1;
		16'hAC67: out_word = 8'hC9;
		16'hAC68: out_word = 8'h3A;
		16'hAC69: out_word = 8'h0D;
		16'hAC6A: out_word = 8'hEC;
		16'hAC6B: out_word = 8'hCB;
		16'hAC6C: out_word = 8'h5F;
		16'hAC6D: out_word = 8'h37;
		16'hAC6E: out_word = 8'hC8;
		16'hAC6F: out_word = 8'hCD;
		16'hAC70: out_word = 8'hB4;
		16'hAC71: out_word = 8'h30;
		16'hAC72: out_word = 8'h21;
		16'hAC73: out_word = 8'h20;
		16'hAC74: out_word = 8'h00;
		16'hAC75: out_word = 8'h19;
		16'hAC76: out_word = 8'hCB;
		16'hAC77: out_word = 8'h5E;
		16'hAC78: out_word = 8'h37;
		16'hAC79: out_word = 8'hC8;
		16'hAC7A: out_word = 8'h18;
		16'hAC7B: out_word = 8'h12;
		16'hAC7C: out_word = 8'h3A;
		16'hAC7D: out_word = 8'h0D;
		16'hAC7E: out_word = 8'hEC;
		16'hAC7F: out_word = 8'hCB;
		16'hAC80: out_word = 8'h5F;
		16'hAC81: out_word = 8'h37;
		16'hAC82: out_word = 8'hC8;
		16'hAC83: out_word = 8'hCD;
		16'hAC84: out_word = 8'hB4;
		16'hAC85: out_word = 8'h30;
		16'hAC86: out_word = 8'h21;
		16'hAC87: out_word = 8'h20;
		16'hAC88: out_word = 8'h00;
		16'hAC89: out_word = 8'h19;
		16'hAC8A: out_word = 8'hCB;
		16'hAC8B: out_word = 8'h46;
		16'hAC8C: out_word = 8'h37;
		16'hAC8D: out_word = 8'hC8;
		16'hAC8E: out_word = 8'h3E;
		16'hAC8F: out_word = 8'h02;
		16'hAC90: out_word = 8'hCD;
		16'hAC91: out_word = 8'hB4;
		16'hAC92: out_word = 8'h30;
		16'hAC93: out_word = 8'h21;
		16'hAC94: out_word = 8'h20;
		16'hAC95: out_word = 8'h00;
		16'hAC96: out_word = 8'h19;
		16'hAC97: out_word = 8'hCB;
		16'hAC98: out_word = 8'h46;
		16'hAC99: out_word = 8'h20;
		16'hAC9A: out_word = 8'h08;
		16'hAC9B: out_word = 8'h0D;
		16'hAC9C: out_word = 8'hF2;
		16'hAC9D: out_word = 8'h90;
		16'hAC9E: out_word = 8'h2C;
		16'hAC9F: out_word = 8'h0E;
		16'hACA0: out_word = 8'h00;
		16'hACA1: out_word = 8'h3E;
		16'hACA2: out_word = 8'h01;
		16'hACA3: out_word = 8'h21;
		16'hACA4: out_word = 8'h00;
		16'hACA5: out_word = 8'hEC;
		16'hACA6: out_word = 8'h11;
		16'hACA7: out_word = 8'h03;
		16'hACA8: out_word = 8'hEC;
		16'hACA9: out_word = 8'hF6;
		16'hACAA: out_word = 8'h80;
		16'hACAB: out_word = 8'h77;
		16'hACAC: out_word = 8'h12;
		16'hACAD: out_word = 8'h23;
		16'hACAE: out_word = 8'h13;
		16'hACAF: out_word = 8'h3E;
		16'hACB0: out_word = 8'h00;
		16'hACB1: out_word = 8'h77;
		16'hACB2: out_word = 8'h12;
		16'hACB3: out_word = 8'h23;
		16'hACB4: out_word = 8'h13;
		16'hACB5: out_word = 8'h79;
		16'hACB6: out_word = 8'h77;
		16'hACB7: out_word = 8'h12;
		16'hACB8: out_word = 8'h21;
		16'hACB9: out_word = 8'h00;
		16'hACBA: out_word = 8'h00;
		16'hACBB: out_word = 8'h22;
		16'hACBC: out_word = 8'h06;
		16'hACBD: out_word = 8'hEC;
		16'hACBE: out_word = 8'hCD;
		16'hACBF: out_word = 8'h5F;
		16'hACC0: out_word = 8'h33;
		16'hACC1: out_word = 8'hCD;
		16'hACC2: out_word = 8'h67;
		16'hACC3: out_word = 8'h3C;
		16'hACC4: out_word = 8'hDD;
		16'hACC5: out_word = 8'hE5;
		16'hACC6: out_word = 8'hCD;
		16'hACC7: out_word = 8'h20;
		16'hACC8: out_word = 8'h1F;
		16'hACC9: out_word = 8'hCD;
		16'hACCA: out_word = 8'h6B;
		16'hACCB: out_word = 8'h02;
		16'hACCC: out_word = 8'hCD;
		16'hACCD: out_word = 8'h45;
		16'hACCE: out_word = 8'h1F;
		16'hACCF: out_word = 8'hDD;
		16'hACD0: out_word = 8'hE1;
		16'hACD1: out_word = 8'h3A;
		16'hACD2: out_word = 8'h3A;
		16'hACD3: out_word = 8'h5C;
		16'hACD4: out_word = 8'h3C;
		16'hACD5: out_word = 8'h20;
		16'hACD6: out_word = 8'h18;
		16'hACD7: out_word = 8'h21;
		16'hACD8: out_word = 8'h0D;
		16'hACD9: out_word = 8'hEC;
		16'hACDA: out_word = 8'hCB;
		16'hACDB: out_word = 8'h9E;
		16'hACDC: out_word = 8'hCD;
		16'hACDD: out_word = 8'h5E;
		16'hACDE: out_word = 8'h36;
		16'hACDF: out_word = 8'h3A;
		16'hACE0: out_word = 8'h0E;
		16'hACE1: out_word = 8'hEC;
		16'hACE2: out_word = 8'hFE;
		16'hACE3: out_word = 8'h04;
		16'hACE4: out_word = 8'hC4;
		16'hACE5: out_word = 8'h2F;
		16'hACE6: out_word = 8'h15;
		16'hACE7: out_word = 8'hCD;
		16'hACE8: out_word = 8'hFA;
		16'hACE9: out_word = 8'h26;
		16'hACEA: out_word = 8'hCD;
		16'hACEB: out_word = 8'h07;
		16'hACEC: out_word = 8'h2A;
		16'hACED: out_word = 8'h37;
		16'hACEE: out_word = 8'hC9;
		16'hACEF: out_word = 8'h21;
		16'hACF0: out_word = 8'h00;
		16'hACF1: out_word = 8'hEC;
		16'hACF2: out_word = 8'h11;
		16'hACF3: out_word = 8'h03;
		16'hACF4: out_word = 8'hEC;
		16'hACF5: out_word = 8'h1A;
		16'hACF6: out_word = 8'hCB;
		16'hACF7: out_word = 8'hBF;
		16'hACF8: out_word = 8'h77;
		16'hACF9: out_word = 8'h23;
		16'hACFA: out_word = 8'h13;
		16'hACFB: out_word = 8'h1A;
		16'hACFC: out_word = 8'h77;
		16'hACFD: out_word = 8'h23;
		16'hACFE: out_word = 8'h13;
		16'hACFF: out_word = 8'h1A;
		16'hAD00: out_word = 8'h77;
		16'hAD01: out_word = 8'hCD;
		16'hAD02: out_word = 8'h63;
		16'hAD03: out_word = 8'h3C;
		16'hAD04: out_word = 8'h38;
		16'hAD05: out_word = 8'h04;
		16'hAD06: out_word = 8'hED;
		16'hAD07: out_word = 8'h4B;
		16'hAD08: out_word = 8'h06;
		16'hAD09: out_word = 8'hEC;
		16'hAD0A: out_word = 8'h2A;
		16'hAD0B: out_word = 8'h06;
		16'hAD0C: out_word = 8'hEC;
		16'hAD0D: out_word = 8'hB7;
		16'hAD0E: out_word = 8'hED;
		16'hAD0F: out_word = 8'h42;
		16'hAD10: out_word = 8'hF5;
		16'hAD11: out_word = 8'hE5;
		16'hAD12: out_word = 8'hCD;
		16'hAD13: out_word = 8'h07;
		16'hAD14: out_word = 8'h2A;
		16'hAD15: out_word = 8'hE1;
		16'hAD16: out_word = 8'hF1;
		16'hAD17: out_word = 8'h38;
		16'hAD18: out_word = 8'h11;
		16'hAD19: out_word = 8'h28;
		16'hAD1A: out_word = 8'h2A;
		16'hAD1B: out_word = 8'hE5;
		16'hAD1C: out_word = 8'h78;
		16'hAD1D: out_word = 8'hCD;
		16'hAD1E: out_word = 8'h5B;
		16'hAD1F: out_word = 8'h2B;
		16'hAD20: out_word = 8'hE1;
		16'hAD21: out_word = 8'h30;
		16'hAD22: out_word = 8'h22;
		16'hAD23: out_word = 8'h2B;
		16'hAD24: out_word = 8'h7C;
		16'hAD25: out_word = 8'hB5;
		16'hAD26: out_word = 8'h20;
		16'hAD27: out_word = 8'hF3;
		16'hAD28: out_word = 8'h18;
		16'hAD29: out_word = 8'h1B;
		16'hAD2A: out_word = 8'hE5;
		16'hAD2B: out_word = 8'h21;
		16'hAD2C: out_word = 8'h0D;
		16'hAD2D: out_word = 8'hEC;
		16'hAD2E: out_word = 8'hCB;
		16'hAD2F: out_word = 8'hBE;
		16'hAD30: out_word = 8'hE1;
		16'hAD31: out_word = 8'hEB;
		16'hAD32: out_word = 8'h21;
		16'hAD33: out_word = 8'h00;
		16'hAD34: out_word = 8'h00;
		16'hAD35: out_word = 8'hB7;
		16'hAD36: out_word = 8'hED;
		16'hAD37: out_word = 8'h52;
		16'hAD38: out_word = 8'hE5;
		16'hAD39: out_word = 8'h78;
		16'hAD3A: out_word = 8'hCD;
		16'hAD3B: out_word = 8'h78;
		16'hAD3C: out_word = 8'h2B;
		16'hAD3D: out_word = 8'hE1;
		16'hAD3E: out_word = 8'h30;
		16'hAD3F: out_word = 8'h05;
		16'hAD40: out_word = 8'h2B;
		16'hAD41: out_word = 8'h7C;
		16'hAD42: out_word = 8'hB5;
		16'hAD43: out_word = 8'h20;
		16'hAD44: out_word = 8'hF3;
		16'hAD45: out_word = 8'h21;
		16'hAD46: out_word = 8'h0D;
		16'hAD47: out_word = 8'hEC;
		16'hAD48: out_word = 8'hCB;
		16'hAD49: out_word = 8'hFE;
		16'hAD4A: out_word = 8'hCD;
		16'hAD4B: out_word = 8'h11;
		16'hAD4C: out_word = 8'h2A;
		16'hAD4D: out_word = 8'h3E;
		16'hAD4E: out_word = 8'h17;
		16'hAD4F: out_word = 8'hCD;
		16'hAD50: out_word = 8'h96;
		16'hAD51: out_word = 8'h3A;
		16'hAD52: out_word = 8'hB7;
		16'hAD53: out_word = 8'hC9;
		16'hAD54: out_word = 8'h21;
		16'hAD55: out_word = 8'h00;
		16'hAD56: out_word = 8'hEC;
		16'hAD57: out_word = 8'hCB;
		16'hAD58: out_word = 8'h7E;
		16'hAD59: out_word = 8'h28;
		16'hAD5A: out_word = 8'h07;
		16'hAD5B: out_word = 8'h2A;
		16'hAD5C: out_word = 8'h06;
		16'hAD5D: out_word = 8'hEC;
		16'hAD5E: out_word = 8'h23;
		16'hAD5F: out_word = 8'h22;
		16'hAD60: out_word = 8'h06;
		16'hAD61: out_word = 8'hEC;
		16'hAD62: out_word = 8'h21;
		16'hAD63: out_word = 8'h00;
		16'hAD64: out_word = 8'hEC;
		16'hAD65: out_word = 8'h7E;
		16'hAD66: out_word = 8'h23;
		16'hAD67: out_word = 8'h46;
		16'hAD68: out_word = 8'h23;
		16'hAD69: out_word = 8'h4E;
		16'hAD6A: out_word = 8'hE5;
		16'hAD6B: out_word = 8'hE6;
		16'hAD6C: out_word = 8'h0F;
		16'hAD6D: out_word = 8'h21;
		16'hAD6E: out_word = 8'h85;
		16'hAD6F: out_word = 8'h2D;
		16'hAD70: out_word = 8'hCD;
		16'hAD71: out_word = 8'hCE;
		16'hAD72: out_word = 8'h3F;
		16'hAD73: out_word = 8'h5D;
		16'hAD74: out_word = 8'hE1;
		16'hAD75: out_word = 8'h28;
		16'hAD76: out_word = 8'h02;
		16'hAD77: out_word = 8'h3E;
		16'hAD78: out_word = 8'h0D;
		16'hAD79: out_word = 8'h71;
		16'hAD7A: out_word = 8'h2B;
		16'hAD7B: out_word = 8'h70;
		16'hAD7C: out_word = 8'h2B;
		16'hAD7D: out_word = 8'hF5;
		16'hAD7E: out_word = 8'h7E;
		16'hAD7F: out_word = 8'hE6;
		16'hAD80: out_word = 8'hF0;
		16'hAD81: out_word = 8'hB3;
		16'hAD82: out_word = 8'h77;
		16'hAD83: out_word = 8'hF1;
		16'hAD84: out_word = 8'hC9;
		16'hAD85: out_word = 8'h03;
		16'hAD86: out_word = 8'h02;
		16'hAD87: out_word = 8'hAC;
		16'hAD88: out_word = 8'h2D;
		16'hAD89: out_word = 8'h04;
		16'hAD8A: out_word = 8'hE9;
		16'hAD8B: out_word = 8'h2D;
		16'hAD8C: out_word = 8'h01;
		16'hAD8D: out_word = 8'h8F;
		16'hAD8E: out_word = 8'h2D;
		16'hAD8F: out_word = 8'hCD;
		16'hAD90: out_word = 8'hB7;
		16'hAD91: out_word = 8'h32;
		16'hAD92: out_word = 8'hCD;
		16'hAD93: out_word = 8'h0E;
		16'hAD94: out_word = 8'h2E;
		16'hAD95: out_word = 8'h30;
		16'hAD96: out_word = 8'h07;
		16'hAD97: out_word = 8'hFE;
		16'hAD98: out_word = 8'h00;
		16'hAD99: out_word = 8'h28;
		16'hAD9A: out_word = 8'hF7;
		16'hAD9B: out_word = 8'h2E;
		16'hAD9C: out_word = 8'h01;
		16'hAD9D: out_word = 8'hC9;
		16'hAD9E: out_word = 8'h0C;
		16'hAD9F: out_word = 8'h06;
		16'hADA0: out_word = 8'h00;
		16'hADA1: out_word = 8'h2A;
		16'hADA2: out_word = 8'hDB;
		16'hADA3: out_word = 8'hF9;
		16'hADA4: out_word = 8'h79;
		16'hADA5: out_word = 8'hBE;
		16'hADA6: out_word = 8'h38;
		16'hADA7: out_word = 8'hE7;
		16'hADA8: out_word = 8'h06;
		16'hADA9: out_word = 8'h00;
		16'hADAA: out_word = 8'h0E;
		16'hADAB: out_word = 8'h00;
		16'hADAC: out_word = 8'hE5;
		16'hADAD: out_word = 8'h21;
		16'hADAE: out_word = 8'hEE;
		16'hADAF: out_word = 8'hF6;
		16'hADB0: out_word = 8'h7E;
		16'hADB1: out_word = 8'hB9;
		16'hADB2: out_word = 8'h20;
		16'hADB3: out_word = 8'h0A;
		16'hADB4: out_word = 8'h23;
		16'hADB5: out_word = 8'h7E;
		16'hADB6: out_word = 8'hB8;
		16'hADB7: out_word = 8'h20;
		16'hADB8: out_word = 8'h05;
		16'hADB9: out_word = 8'h21;
		16'hADBA: out_word = 8'h00;
		16'hADBB: out_word = 8'hEC;
		16'hADBC: out_word = 8'hCB;
		16'hADBD: out_word = 8'hBE;
		16'hADBE: out_word = 8'hE1;
		16'hADBF: out_word = 8'hCD;
		16'hADC0: out_word = 8'hB4;
		16'hADC1: out_word = 8'h30;
		16'hADC2: out_word = 8'hCD;
		16'hADC3: out_word = 8'h0E;
		16'hADC4: out_word = 8'h2E;
		16'hADC5: out_word = 8'h30;
		16'hADC6: out_word = 8'h07;
		16'hADC7: out_word = 8'hFE;
		16'hADC8: out_word = 8'h00;
		16'hADC9: out_word = 8'h28;
		16'hADCA: out_word = 8'hE1;
		16'hADCB: out_word = 8'h2E;
		16'hADCC: out_word = 8'h02;
		16'hADCD: out_word = 8'hC9;
		16'hADCE: out_word = 8'h21;
		16'hADCF: out_word = 8'h20;
		16'hADD0: out_word = 8'h00;
		16'hADD1: out_word = 8'h19;
		16'hADD2: out_word = 8'hCB;
		16'hADD3: out_word = 8'h5E;
		16'hADD4: out_word = 8'h28;
		16'hADD5: out_word = 8'h05;
		16'hADD6: out_word = 8'h2E;
		16'hADD7: out_word = 8'h08;
		16'hADD8: out_word = 8'h3E;
		16'hADD9: out_word = 8'h0D;
		16'hADDA: out_word = 8'hC9;
		16'hADDB: out_word = 8'h21;
		16'hADDC: out_word = 8'hF3;
		16'hADDD: out_word = 8'hF6;
		16'hADDE: out_word = 8'h0C;
		16'hADDF: out_word = 8'h7E;
		16'hADE0: out_word = 8'hB9;
		16'hADE1: out_word = 8'h06;
		16'hADE2: out_word = 8'h00;
		16'hADE3: out_word = 8'h30;
		16'hADE4: out_word = 8'hDA;
		16'hADE5: out_word = 8'h06;
		16'hADE6: out_word = 8'h00;
		16'hADE7: out_word = 8'h0E;
		16'hADE8: out_word = 8'h01;
		16'hADE9: out_word = 8'hCD;
		16'hADEA: out_word = 8'hC3;
		16'hADEB: out_word = 8'h31;
		16'hADEC: out_word = 8'hCD;
		16'hADED: out_word = 8'h0E;
		16'hADEE: out_word = 8'h2E;
		16'hADEF: out_word = 8'h30;
		16'hADF0: out_word = 8'h07;
		16'hADF1: out_word = 8'hFE;
		16'hADF2: out_word = 8'h00;
		16'hADF3: out_word = 8'h28;
		16'hADF4: out_word = 8'hF7;
		16'hADF5: out_word = 8'h2E;
		16'hADF6: out_word = 8'h04;
		16'hADF7: out_word = 8'hC9;
		16'hADF8: out_word = 8'h21;
		16'hADF9: out_word = 8'h20;
		16'hADFA: out_word = 8'h00;
		16'hADFB: out_word = 8'h19;
		16'hADFC: out_word = 8'hCB;
		16'hADFD: out_word = 8'h5E;
		16'hADFE: out_word = 8'h20;
		16'hADFF: out_word = 8'h09;
		16'hAE00: out_word = 8'h0C;
		16'hAE01: out_word = 8'h06;
		16'hAE02: out_word = 8'h00;
		16'hAE03: out_word = 8'h3A;
		16'hAE04: out_word = 8'hF5;
		16'hAE05: out_word = 8'hF6;
		16'hAE06: out_word = 8'hB9;
		16'hAE07: out_word = 8'h30;
		16'hAE08: out_word = 8'hE0;
		16'hAE09: out_word = 8'h2E;
		16'hAE0A: out_word = 8'h08;
		16'hAE0B: out_word = 8'h3E;
		16'hAE0C: out_word = 8'h0D;
		16'hAE0D: out_word = 8'hC9;
		16'hAE0E: out_word = 8'h3E;
		16'hAE0F: out_word = 8'h1F;
		16'hAE10: out_word = 8'hB8;
		16'hAE11: out_word = 8'h3F;
		16'hAE12: out_word = 8'hD0;
		16'hAE13: out_word = 8'h68;
		16'hAE14: out_word = 8'h26;
		16'hAE15: out_word = 8'h00;
		16'hAE16: out_word = 8'h19;
		16'hAE17: out_word = 8'h7E;
		16'hAE18: out_word = 8'h04;
		16'hAE19: out_word = 8'h37;
		16'hAE1A: out_word = 8'hC9;
		16'hAE1B: out_word = 8'h01;
		16'hAE1C: out_word = 8'h14;
		16'hAE1D: out_word = 8'h01;
		16'hAE1E: out_word = 8'h01;
		16'hAE1F: out_word = 8'h21;
		16'hAE20: out_word = 8'h3C;
		16'hAE21: out_word = 8'h5C;
		16'hAE22: out_word = 8'hCB;
		16'hAE23: out_word = 8'h86;
		16'hAE24: out_word = 8'h21;
		16'hAE25: out_word = 8'h1B;
		16'hAE26: out_word = 8'h2E;
		16'hAE27: out_word = 8'h11;
		16'hAE28: out_word = 8'h15;
		16'hAE29: out_word = 8'hEC;
		16'hAE2A: out_word = 8'hC3;
		16'hAE2B: out_word = 8'hBA;
		16'hAE2C: out_word = 8'h3F;
		16'hAE2D: out_word = 8'h21;
		16'hAE2E: out_word = 8'h3C;
		16'hAE2F: out_word = 8'h5C;
		16'hAE30: out_word = 8'hCB;
		16'hAE31: out_word = 8'hC6;
		16'hAE32: out_word = 8'h01;
		16'hAE33: out_word = 8'h00;
		16'hAE34: out_word = 8'h00;
		16'hAE35: out_word = 8'hCD;
		16'hAE36: out_word = 8'h2B;
		16'hAE37: out_word = 8'h37;
		16'hAE38: out_word = 8'h21;
		16'hAE39: out_word = 8'h1D;
		16'hAE3A: out_word = 8'h2E;
		16'hAE3B: out_word = 8'h11;
		16'hAE3C: out_word = 8'h15;
		16'hAE3D: out_word = 8'hEC;
		16'hAE3E: out_word = 8'hC3;
		16'hAE3F: out_word = 8'hBA;
		16'hAE40: out_word = 8'h3F;
		16'hAE41: out_word = 8'h26;
		16'hAE42: out_word = 8'h00;
		16'hAE43: out_word = 8'h68;
		16'hAE44: out_word = 8'h19;
		16'hAE45: out_word = 8'h7E;
		16'hAE46: out_word = 8'hFE;
		16'hAE47: out_word = 8'h00;
		16'hAE48: out_word = 8'h37;
		16'hAE49: out_word = 8'hC0;
		16'hAE4A: out_word = 8'h78;
		16'hAE4B: out_word = 8'hB7;
		16'hAE4C: out_word = 8'h28;
		16'hAE4D: out_word = 8'h0D;
		16'hAE4E: out_word = 8'hE5;
		16'hAE4F: out_word = 8'h2B;
		16'hAE50: out_word = 8'h7E;
		16'hAE51: out_word = 8'hFE;
		16'hAE52: out_word = 8'h00;
		16'hAE53: out_word = 8'h37;
		16'hAE54: out_word = 8'hE1;
		16'hAE55: out_word = 8'hC0;
		16'hAE56: out_word = 8'h7E;
		16'hAE57: out_word = 8'hFE;
		16'hAE58: out_word = 8'h00;
		16'hAE59: out_word = 8'h37;
		16'hAE5A: out_word = 8'hC0;
		16'hAE5B: out_word = 8'h23;
		16'hAE5C: out_word = 8'h04;
		16'hAE5D: out_word = 8'h78;
		16'hAE5E: out_word = 8'hFE;
		16'hAE5F: out_word = 8'h1F;
		16'hAE60: out_word = 8'h38;
		16'hAE61: out_word = 8'hF4;
		16'hAE62: out_word = 8'hC9;
		16'hAE63: out_word = 8'h26;
		16'hAE64: out_word = 8'h00;
		16'hAE65: out_word = 8'h68;
		16'hAE66: out_word = 8'h19;
		16'hAE67: out_word = 8'h7E;
		16'hAE68: out_word = 8'hFE;
		16'hAE69: out_word = 8'h00;
		16'hAE6A: out_word = 8'h37;
		16'hAE6B: out_word = 8'hC0;
		16'hAE6C: out_word = 8'h7E;
		16'hAE6D: out_word = 8'hFE;
		16'hAE6E: out_word = 8'h00;
		16'hAE6F: out_word = 8'h20;
		16'hAE70: out_word = 8'h07;
		16'hAE71: out_word = 8'h78;
		16'hAE72: out_word = 8'hB7;
		16'hAE73: out_word = 8'hC8;
		16'hAE74: out_word = 8'h2B;
		16'hAE75: out_word = 8'h05;
		16'hAE76: out_word = 8'h18;
		16'hAE77: out_word = 8'hF4;
		16'hAE78: out_word = 8'h04;
		16'hAE79: out_word = 8'h37;
		16'hAE7A: out_word = 8'hC9;
		16'hAE7B: out_word = 8'h26;
		16'hAE7C: out_word = 8'h00;
		16'hAE7D: out_word = 8'h68;
		16'hAE7E: out_word = 8'h19;
		16'hAE7F: out_word = 8'h7E;
		16'hAE80: out_word = 8'hC9;
		16'hAE81: out_word = 8'h21;
		16'hAE82: out_word = 8'h0D;
		16'hAE83: out_word = 8'hEC;
		16'hAE84: out_word = 8'hB7;
		16'hAE85: out_word = 8'hCB;
		16'hAE86: out_word = 8'h46;
		16'hAE87: out_word = 8'hC0;
		16'hAE88: out_word = 8'hC5;
		16'hAE89: out_word = 8'hF5;
		16'hAE8A: out_word = 8'hCD;
		16'hAE8B: out_word = 8'hB4;
		16'hAE8C: out_word = 8'h30;
		16'hAE8D: out_word = 8'hF1;
		16'hAE8E: out_word = 8'hCD;
		16'hAE8F: out_word = 8'hAC;
		16'hAE90: out_word = 8'h16;
		16'hAE91: out_word = 8'hF5;
		16'hAE92: out_word = 8'hEB;
		16'hAE93: out_word = 8'hCD;
		16'hAE94: out_word = 8'h04;
		16'hAE95: out_word = 8'h36;
		16'hAE96: out_word = 8'hEB;
		16'hAE97: out_word = 8'hF1;
		16'hAE98: out_word = 8'h3F;
		16'hAE99: out_word = 8'h28;
		16'hAE9A: out_word = 8'h31;
		16'hAE9B: out_word = 8'hF5;
		16'hAE9C: out_word = 8'h06;
		16'hAE9D: out_word = 8'h00;
		16'hAE9E: out_word = 8'h0C;
		16'hAE9F: out_word = 8'h3A;
		16'hAEA0: out_word = 8'h15;
		16'hAEA1: out_word = 8'hEC;
		16'hAEA2: out_word = 8'hB9;
		16'hAEA3: out_word = 8'h38;
		16'hAEA4: out_word = 8'h23;
		16'hAEA5: out_word = 8'h7E;
		16'hAEA6: out_word = 8'h5F;
		16'hAEA7: out_word = 8'hE6;
		16'hAEA8: out_word = 8'hD7;
		16'hAEA9: out_word = 8'hBE;
		16'hAEAA: out_word = 8'h77;
		16'hAEAB: out_word = 8'h7B;
		16'hAEAC: out_word = 8'hCB;
		16'hAEAD: out_word = 8'hCE;
		16'hAEAE: out_word = 8'hF5;
		16'hAEAF: out_word = 8'hCD;
		16'hAEB0: out_word = 8'hB4;
		16'hAEB1: out_word = 8'h30;
		16'hAEB2: out_word = 8'hF1;
		16'hAEB3: out_word = 8'h28;
		16'hAEB4: out_word = 8'h0D;
		16'hAEB5: out_word = 8'hCB;
		16'hAEB6: out_word = 8'h87;
		16'hAEB7: out_word = 8'hCD;
		16'hAEB8: out_word = 8'hD3;
		16'hAEB9: out_word = 8'h2E;
		16'hAEBA: out_word = 8'h30;
		16'hAEBB: out_word = 8'h10;
		16'hAEBC: out_word = 8'hCD;
		16'hAEBD: out_word = 8'hF4;
		16'hAEBE: out_word = 8'h35;
		16'hAEBF: out_word = 8'hF1;
		16'hAEC0: out_word = 8'h18;
		16'hAEC1: out_word = 8'hCC;
		16'hAEC2: out_word = 8'hCD;
		16'hAEC3: out_word = 8'h41;
		16'hAEC4: out_word = 8'h2E;
		16'hAEC5: out_word = 8'hF1;
		16'hAEC6: out_word = 8'h18;
		16'hAEC7: out_word = 8'hC6;
		16'hAEC8: out_word = 8'hF1;
		16'hAEC9: out_word = 8'hCD;
		16'hAECA: out_word = 8'h6E;
		16'hAECB: out_word = 8'h31;
		16'hAECC: out_word = 8'hC1;
		16'hAECD: out_word = 8'hC9;
		16'hAECE: out_word = 8'hCD;
		16'hAECF: out_word = 8'hB4;
		16'hAED0: out_word = 8'h30;
		16'hAED1: out_word = 8'h3E;
		16'hAED2: out_word = 8'h09;
		16'hAED3: out_word = 8'hC5;
		16'hAED4: out_word = 8'hD5;
		16'hAED5: out_word = 8'h41;
		16'hAED6: out_word = 8'h21;
		16'hAED7: out_word = 8'hEF;
		16'hAED8: out_word = 8'h2E;
		16'hAED9: out_word = 8'h4F;
		16'hAEDA: out_word = 8'hC5;
		16'hAEDB: out_word = 8'hCD;
		16'hAEDC: out_word = 8'h75;
		16'hAEDD: out_word = 8'h16;
		16'hAEDE: out_word = 8'hC1;
		16'hAEDF: out_word = 8'h79;
		16'hAEE0: out_word = 8'h30;
		16'hAEE1: out_word = 8'h0A;
		16'hAEE2: out_word = 8'h48;
		16'hAEE3: out_word = 8'hCD;
		16'hAEE4: out_word = 8'hB4;
		16'hAEE5: out_word = 8'h30;
		16'hAEE6: out_word = 8'h21;
		16'hAEE7: out_word = 8'h20;
		16'hAEE8: out_word = 8'h00;
		16'hAEE9: out_word = 8'h19;
		16'hAEEA: out_word = 8'h77;
		16'hAEEB: out_word = 8'h37;
		16'hAEEC: out_word = 8'hD1;
		16'hAEED: out_word = 8'hC1;
		16'hAEEE: out_word = 8'hC9;
		16'hAEEF: out_word = 8'h00;
		16'hAEF0: out_word = 8'h00;
		16'hAEF1: out_word = 8'h00;
		16'hAEF2: out_word = 8'h00;
		16'hAEF3: out_word = 8'h00;
		16'hAEF4: out_word = 8'h00;
		16'hAEF5: out_word = 8'h00;
		16'hAEF6: out_word = 8'h00;
		16'hAEF7: out_word = 8'h00;
		16'hAEF8: out_word = 8'h00;
		16'hAEF9: out_word = 8'h00;
		16'hAEFA: out_word = 8'h00;
		16'hAEFB: out_word = 8'h00;
		16'hAEFC: out_word = 8'h00;
		16'hAEFD: out_word = 8'h00;
		16'hAEFE: out_word = 8'h00;
		16'hAEFF: out_word = 8'h00;
		16'hAF00: out_word = 8'h00;
		16'hAF01: out_word = 8'h00;
		16'hAF02: out_word = 8'h00;
		16'hAF03: out_word = 8'h00;
		16'hAF04: out_word = 8'h00;
		16'hAF05: out_word = 8'h00;
		16'hAF06: out_word = 8'h00;
		16'hAF07: out_word = 8'h00;
		16'hAF08: out_word = 8'h00;
		16'hAF09: out_word = 8'h00;
		16'hAF0A: out_word = 8'h00;
		16'hAF0B: out_word = 8'h00;
		16'hAF0C: out_word = 8'h00;
		16'hAF0D: out_word = 8'h00;
		16'hAF0E: out_word = 8'h00;
		16'hAF0F: out_word = 8'h09;
		16'hAF10: out_word = 8'h00;
		16'hAF11: out_word = 8'h00;
		16'hAF12: out_word = 8'hC5;
		16'hAF13: out_word = 8'hCD;
		16'hAF14: out_word = 8'hB4;
		16'hAF15: out_word = 8'h30;
		16'hAF16: out_word = 8'hC5;
		16'hAF17: out_word = 8'h21;
		16'hAF18: out_word = 8'h20;
		16'hAF19: out_word = 8'h00;
		16'hAF1A: out_word = 8'h19;
		16'hAF1B: out_word = 8'hCB;
		16'hAF1C: out_word = 8'h4E;
		16'hAF1D: out_word = 8'h3E;
		16'hAF1E: out_word = 8'h00;
		16'hAF1F: out_word = 8'h28;
		16'hAF20: out_word = 8'h10;
		16'hAF21: out_word = 8'h0C;
		16'hAF22: out_word = 8'h21;
		16'hAF23: out_word = 8'h23;
		16'hAF24: out_word = 8'h00;
		16'hAF25: out_word = 8'h19;
		16'hAF26: out_word = 8'hEB;
		16'hAF27: out_word = 8'h3A;
		16'hAF28: out_word = 8'h15;
		16'hAF29: out_word = 8'hEC;
		16'hAF2A: out_word = 8'hB9;
		16'hAF2B: out_word = 8'h30;
		16'hAF2C: out_word = 8'hEA;
		16'hAF2D: out_word = 8'h0D;
		16'hAF2E: out_word = 8'hCD;
		16'hAF2F: out_word = 8'hC9;
		16'hAF30: out_word = 8'h31;
		16'hAF31: out_word = 8'hE1;
		16'hAF32: out_word = 8'hE5;
		16'hAF33: out_word = 8'hCD;
		16'hAF34: out_word = 8'hB4;
		16'hAF35: out_word = 8'h30;
		16'hAF36: out_word = 8'hE1;
		16'hAF37: out_word = 8'h47;
		16'hAF38: out_word = 8'h79;
		16'hAF39: out_word = 8'hBD;
		16'hAF3A: out_word = 8'h78;
		16'hAF3B: out_word = 8'hF5;
		16'hAF3C: out_word = 8'h20;
		16'hAF3D: out_word = 8'h03;
		16'hAF3E: out_word = 8'h44;
		16'hAF3F: out_word = 8'h18;
		16'hAF40: out_word = 8'h09;
		16'hAF41: out_word = 8'hF5;
		16'hAF42: out_word = 8'hE5;
		16'hAF43: out_word = 8'h06;
		16'hAF44: out_word = 8'h00;
		16'hAF45: out_word = 8'hCD;
		16'hAF46: out_word = 8'h41;
		16'hAF47: out_word = 8'h2E;
		16'hAF48: out_word = 8'hE1;
		16'hAF49: out_word = 8'hF1;
		16'hAF4A: out_word = 8'hE5;
		16'hAF4B: out_word = 8'h21;
		16'hAF4C: out_word = 8'hF4;
		16'hAF4D: out_word = 8'hF6;
		16'hAF4E: out_word = 8'hCB;
		16'hAF4F: out_word = 8'hC6;
		16'hAF50: out_word = 8'h28;
		16'hAF51: out_word = 8'h02;
		16'hAF52: out_word = 8'hCB;
		16'hAF53: out_word = 8'h86;
		16'hAF54: out_word = 8'hCD;
		16'hAF55: out_word = 8'hC1;
		16'hAF56: out_word = 8'h16;
		16'hAF57: out_word = 8'hF5;
		16'hAF58: out_word = 8'hC5;
		16'hAF59: out_word = 8'hD5;
		16'hAF5A: out_word = 8'h21;
		16'hAF5B: out_word = 8'hF4;
		16'hAF5C: out_word = 8'hF6;
		16'hAF5D: out_word = 8'hCB;
		16'hAF5E: out_word = 8'h46;
		16'hAF5F: out_word = 8'h20;
		16'hAF60: out_word = 8'h0E;
		16'hAF61: out_word = 8'h06;
		16'hAF62: out_word = 8'h00;
		16'hAF63: out_word = 8'hCD;
		16'hAF64: out_word = 8'hD4;
		16'hAF65: out_word = 8'h2B;
		16'hAF66: out_word = 8'h38;
		16'hAF67: out_word = 8'h07;
		16'hAF68: out_word = 8'hCD;
		16'hAF69: out_word = 8'h80;
		16'hAF6A: out_word = 8'h2F;
		16'hAF6B: out_word = 8'hD1;
		16'hAF6C: out_word = 8'hC1;
		16'hAF6D: out_word = 8'h18;
		16'hAF6E: out_word = 8'h05;
		16'hAF6F: out_word = 8'hE1;
		16'hAF70: out_word = 8'hC1;
		16'hAF71: out_word = 8'hCD;
		16'hAF72: out_word = 8'h04;
		16'hAF73: out_word = 8'h36;
		16'hAF74: out_word = 8'hF1;
		16'hAF75: out_word = 8'h0D;
		16'hAF76: out_word = 8'h47;
		16'hAF77: out_word = 8'hE1;
		16'hAF78: out_word = 8'hF1;
		16'hAF79: out_word = 8'h78;
		16'hAF7A: out_word = 8'hC2;
		16'hAF7B: out_word = 8'h32;
		16'hAF7C: out_word = 8'h2F;
		16'hAF7D: out_word = 8'h37;
		16'hAF7E: out_word = 8'hC1;
		16'hAF7F: out_word = 8'hC9;
		16'hAF80: out_word = 8'h21;
		16'hAF81: out_word = 8'h20;
		16'hAF82: out_word = 8'h00;
		16'hAF83: out_word = 8'h19;
		16'hAF84: out_word = 8'h7E;
		16'hAF85: out_word = 8'hCB;
		16'hAF86: out_word = 8'h46;
		16'hAF87: out_word = 8'h20;
		16'hAF88: out_word = 8'h29;
		16'hAF89: out_word = 8'hF5;
		16'hAF8A: out_word = 8'hC5;
		16'hAF8B: out_word = 8'h79;
		16'hAF8C: out_word = 8'hB7;
		16'hAF8D: out_word = 8'h20;
		16'hAF8E: out_word = 8'h15;
		16'hAF8F: out_word = 8'hC5;
		16'hAF90: out_word = 8'h2A;
		16'hAF91: out_word = 8'h9A;
		16'hAF92: out_word = 8'hFC;
		16'hAF93: out_word = 8'hCD;
		16'hAF94: out_word = 8'h4A;
		16'hAF95: out_word = 8'h33;
		16'hAF96: out_word = 8'h22;
		16'hAF97: out_word = 8'h9A;
		16'hAF98: out_word = 8'hFC;
		16'hAF99: out_word = 8'h3A;
		16'hAF9A: out_word = 8'hDB;
		16'hAF9B: out_word = 8'hF9;
		16'hAF9C: out_word = 8'h4F;
		16'hAF9D: out_word = 8'h0D;
		16'hAF9E: out_word = 8'hCD;
		16'hAF9F: out_word = 8'hB7;
		16'hAFA0: out_word = 8'h32;
		16'hAFA1: out_word = 8'hC1;
		16'hAFA2: out_word = 8'h18;
		16'hAFA3: out_word = 8'h04;
		16'hAFA4: out_word = 8'h0D;
		16'hAFA5: out_word = 8'hCD;
		16'hAFA6: out_word = 8'hB4;
		16'hAFA7: out_word = 8'h30;
		16'hAFA8: out_word = 8'hC1;
		16'hAFA9: out_word = 8'hF1;
		16'hAFAA: out_word = 8'h21;
		16'hAFAB: out_word = 8'h20;
		16'hAFAC: out_word = 8'h00;
		16'hAFAD: out_word = 8'h19;
		16'hAFAE: out_word = 8'hCB;
		16'hAFAF: out_word = 8'h8E;
		16'hAFB0: out_word = 8'hB6;
		16'hAFB1: out_word = 8'h77;
		16'hAFB2: out_word = 8'h41;
		16'hAFB3: out_word = 8'hCD;
		16'hAFB4: out_word = 8'hB4;
		16'hAFB5: out_word = 8'h30;
		16'hAFB6: out_word = 8'hCD;
		16'hAFB7: out_word = 8'hDF;
		16'hAFB8: out_word = 8'h30;
		16'hAFB9: out_word = 8'hC3;
		16'hAFBA: out_word = 8'h48;
		16'hAFBB: out_word = 8'h16;
		16'hAFBC: out_word = 8'hCD;
		16'hAFBD: out_word = 8'h84;
		16'hAFBE: out_word = 8'h30;
		16'hAFBF: out_word = 8'hE5;
		16'hAFC0: out_word = 8'hCD;
		16'hAFC1: out_word = 8'h95;
		16'hAFC2: out_word = 8'h30;
		16'hAFC3: out_word = 8'h28;
		16'hAFC4: out_word = 8'h32;
		16'hAFC5: out_word = 8'hCD;
		16'hAFC6: out_word = 8'h5B;
		16'hAFC7: out_word = 8'h2B;
		16'hAFC8: out_word = 8'hE1;
		16'hAFC9: out_word = 8'h30;
		16'hAFCA: out_word = 8'h2D;
		16'hAFCB: out_word = 8'hCD;
		16'hAFCC: out_word = 8'h1A;
		16'hAFCD: out_word = 8'h2A;
		16'hAFCE: out_word = 8'hF5;
		16'hAFCF: out_word = 8'hE5;
		16'hAFD0: out_word = 8'hCD;
		16'hAFD1: out_word = 8'h12;
		16'hAFD2: out_word = 8'h2F;
		16'hAFD3: out_word = 8'hE1;
		16'hAFD4: out_word = 8'hF1;
		16'hAFD5: out_word = 8'hFE;
		16'hAFD6: out_word = 8'h20;
		16'hAFD7: out_word = 8'h28;
		16'hAFD8: out_word = 8'hE6;
		16'hAFD9: out_word = 8'hE5;
		16'hAFDA: out_word = 8'hCD;
		16'hAFDB: out_word = 8'h95;
		16'hAFDC: out_word = 8'h30;
		16'hAFDD: out_word = 8'h28;
		16'hAFDE: out_word = 8'h18;
		16'hAFDF: out_word = 8'hCD;
		16'hAFE0: out_word = 8'h5B;
		16'hAFE1: out_word = 8'h2B;
		16'hAFE2: out_word = 8'hE1;
		16'hAFE3: out_word = 8'h30;
		16'hAFE4: out_word = 8'h13;
		16'hAFE5: out_word = 8'hCD;
		16'hAFE6: out_word = 8'h1A;
		16'hAFE7: out_word = 8'h2A;
		16'hAFE8: out_word = 8'hFE;
		16'hAFE9: out_word = 8'h20;
		16'hAFEA: out_word = 8'h28;
		16'hAFEB: out_word = 8'h07;
		16'hAFEC: out_word = 8'hE5;
		16'hAFED: out_word = 8'hCD;
		16'hAFEE: out_word = 8'h12;
		16'hAFEF: out_word = 8'h2F;
		16'hAFF0: out_word = 8'hE1;
		16'hAFF1: out_word = 8'h18;
		16'hAFF2: out_word = 8'hE6;
		16'hAFF3: out_word = 8'hE5;
		16'hAFF4: out_word = 8'hCD;
		16'hAFF5: out_word = 8'h78;
		16'hAFF6: out_word = 8'h2B;
		16'hAFF7: out_word = 8'hE1;
		16'hAFF8: out_word = 8'h78;
		16'hAFF9: out_word = 8'hF5;
		16'hAFFA: out_word = 8'hE5;
		16'hAFFB: out_word = 8'h21;
		16'hAFFC: out_word = 8'hF5;
		16'hAFFD: out_word = 8'hEE;
		16'hAFFE: out_word = 8'hCB;
		16'hAFFF: out_word = 8'h96;
		16'hB000: out_word = 8'h3A;
		16'hB001: out_word = 8'h15;
		16'hB002: out_word = 8'hEC;
		16'hB003: out_word = 8'hC5;
		16'hB004: out_word = 8'h06;
		16'hB005: out_word = 8'h00;
		16'hB006: out_word = 8'h4F;
		16'hB007: out_word = 8'hBF;
		16'hB008: out_word = 8'hCD;
		16'hB009: out_word = 8'h05;
		16'hB00A: out_word = 8'h16;
		16'hB00B: out_word = 8'hC1;
		16'hB00C: out_word = 8'h21;
		16'hB00D: out_word = 8'h0D;
		16'hB00E: out_word = 8'hEC;
		16'hB00F: out_word = 8'hCB;
		16'hB010: out_word = 8'hDE;
		16'hB011: out_word = 8'hE1;
		16'hB012: out_word = 8'hCD;
		16'hB013: out_word = 8'hF8;
		16'hB014: out_word = 8'h29;
		16'hB015: out_word = 8'hF1;
		16'hB016: out_word = 8'hC9;
		16'hB017: out_word = 8'hCD;
		16'hB018: out_word = 8'h84;
		16'hB019: out_word = 8'h30;
		16'hB01A: out_word = 8'hE5;
		16'hB01B: out_word = 8'hCD;
		16'hB01C: out_word = 8'h1A;
		16'hB01D: out_word = 8'h2A;
		16'hB01E: out_word = 8'hE1;
		16'hB01F: out_word = 8'hFE;
		16'hB020: out_word = 8'h00;
		16'hB021: out_word = 8'h37;
		16'hB022: out_word = 8'h28;
		16'hB023: out_word = 8'hD4;
		16'hB024: out_word = 8'hF5;
		16'hB025: out_word = 8'hE5;
		16'hB026: out_word = 8'hCD;
		16'hB027: out_word = 8'h12;
		16'hB028: out_word = 8'h2F;
		16'hB029: out_word = 8'hE1;
		16'hB02A: out_word = 8'hF1;
		16'hB02B: out_word = 8'hFE;
		16'hB02C: out_word = 8'h20;
		16'hB02D: out_word = 8'h20;
		16'hB02E: out_word = 8'hEB;
		16'hB02F: out_word = 8'hCD;
		16'hB030: out_word = 8'h1A;
		16'hB031: out_word = 8'h2A;
		16'hB032: out_word = 8'hFE;
		16'hB033: out_word = 8'h20;
		16'hB034: out_word = 8'h37;
		16'hB035: out_word = 8'h20;
		16'hB036: out_word = 8'hC1;
		16'hB037: out_word = 8'hE5;
		16'hB038: out_word = 8'hCD;
		16'hB039: out_word = 8'h12;
		16'hB03A: out_word = 8'h2F;
		16'hB03B: out_word = 8'hE1;
		16'hB03C: out_word = 8'h18;
		16'hB03D: out_word = 8'hF1;
		16'hB03E: out_word = 8'hCD;
		16'hB03F: out_word = 8'h84;
		16'hB040: out_word = 8'h30;
		16'hB041: out_word = 8'hE5;
		16'hB042: out_word = 8'hCD;
		16'hB043: out_word = 8'hB4;
		16'hB044: out_word = 8'h30;
		16'hB045: out_word = 8'h21;
		16'hB046: out_word = 8'h20;
		16'hB047: out_word = 8'h00;
		16'hB048: out_word = 8'h19;
		16'hB049: out_word = 8'hCB;
		16'hB04A: out_word = 8'h46;
		16'hB04B: out_word = 8'h20;
		16'hB04C: out_word = 8'h0C;
		16'hB04D: out_word = 8'hCD;
		16'hB04E: out_word = 8'h5B;
		16'hB04F: out_word = 8'h2B;
		16'hB050: out_word = 8'h30;
		16'hB051: out_word = 8'h1B;
		16'hB052: out_word = 8'hCD;
		16'hB053: out_word = 8'h12;
		16'hB054: out_word = 8'h2F;
		16'hB055: out_word = 8'hE1;
		16'hB056: out_word = 8'h18;
		16'hB057: out_word = 8'hE9;
		16'hB058: out_word = 8'hE5;
		16'hB059: out_word = 8'h78;
		16'hB05A: out_word = 8'hFE;
		16'hB05B: out_word = 8'h00;
		16'hB05C: out_word = 8'h28;
		16'hB05D: out_word = 8'h0F;
		16'hB05E: out_word = 8'h05;
		16'hB05F: out_word = 8'hCD;
		16'hB060: out_word = 8'h1A;
		16'hB061: out_word = 8'h2A;
		16'hB062: out_word = 8'h04;
		16'hB063: out_word = 8'hFE;
		16'hB064: out_word = 8'h00;
		16'hB065: out_word = 8'h28;
		16'hB066: out_word = 8'h06;
		16'hB067: out_word = 8'h05;
		16'hB068: out_word = 8'hCD;
		16'hB069: out_word = 8'h12;
		16'hB06A: out_word = 8'h2F;
		16'hB06B: out_word = 8'h18;
		16'hB06C: out_word = 8'hEC;
		16'hB06D: out_word = 8'hE1;
		16'hB06E: out_word = 8'h37;
		16'hB06F: out_word = 8'hC3;
		16'hB070: out_word = 8'hF8;
		16'hB071: out_word = 8'h2F;
		16'hB072: out_word = 8'hCD;
		16'hB073: out_word = 8'h84;
		16'hB074: out_word = 8'h30;
		16'hB075: out_word = 8'hCD;
		16'hB076: out_word = 8'h1A;
		16'hB077: out_word = 8'h2A;
		16'hB078: out_word = 8'hFE;
		16'hB079: out_word = 8'h00;
		16'hB07A: out_word = 8'h37;
		16'hB07B: out_word = 8'h28;
		16'hB07C: out_word = 8'hF1;
		16'hB07D: out_word = 8'hE5;
		16'hB07E: out_word = 8'hCD;
		16'hB07F: out_word = 8'h12;
		16'hB080: out_word = 8'h2F;
		16'hB081: out_word = 8'hE1;
		16'hB082: out_word = 8'h18;
		16'hB083: out_word = 8'hF1;
		16'hB084: out_word = 8'h21;
		16'hB085: out_word = 8'h0D;
		16'hB086: out_word = 8'hEC;
		16'hB087: out_word = 8'hCB;
		16'hB088: out_word = 8'h86;
		16'hB089: out_word = 8'hCD;
		16'hB08A: out_word = 8'hEC;
		16'hB08B: out_word = 8'h29;
		16'hB08C: out_word = 8'h21;
		16'hB08D: out_word = 8'hF5;
		16'hB08E: out_word = 8'hEE;
		16'hB08F: out_word = 8'hCB;
		16'hB090: out_word = 8'hD6;
		16'hB091: out_word = 8'h21;
		16'hB092: out_word = 8'hF1;
		16'hB093: out_word = 8'hF6;
		16'hB094: out_word = 8'hC9;
		16'hB095: out_word = 8'hCD;
		16'hB096: out_word = 8'hB4;
		16'hB097: out_word = 8'h30;
		16'hB098: out_word = 8'h21;
		16'hB099: out_word = 8'h20;
		16'hB09A: out_word = 8'h00;
		16'hB09B: out_word = 8'h19;
		16'hB09C: out_word = 8'hCB;
		16'hB09D: out_word = 8'h46;
		16'hB09E: out_word = 8'h28;
		16'hB09F: out_word = 8'h0E;
		16'hB0A0: out_word = 8'h78;
		16'hB0A1: out_word = 8'hFE;
		16'hB0A2: out_word = 8'h00;
		16'hB0A3: out_word = 8'h28;
		16'hB0A4: out_word = 8'h0D;
		16'hB0A5: out_word = 8'h05;
		16'hB0A6: out_word = 8'hCD;
		16'hB0A7: out_word = 8'h1A;
		16'hB0A8: out_word = 8'h2A;
		16'hB0A9: out_word = 8'h04;
		16'hB0AA: out_word = 8'hFE;
		16'hB0AB: out_word = 8'h00;
		16'hB0AC: out_word = 8'h28;
		16'hB0AD: out_word = 8'h04;
		16'hB0AE: out_word = 8'h3E;
		16'hB0AF: out_word = 8'h01;
		16'hB0B0: out_word = 8'hB7;
		16'hB0B1: out_word = 8'hC9;
		16'hB0B2: out_word = 8'hAF;
		16'hB0B3: out_word = 8'hC9;
		16'hB0B4: out_word = 8'h21;
		16'hB0B5: out_word = 8'h16;
		16'hB0B6: out_word = 8'hEC;
		16'hB0B7: out_word = 8'hF5;
		16'hB0B8: out_word = 8'h79;
		16'hB0B9: out_word = 8'h11;
		16'hB0BA: out_word = 8'h23;
		16'hB0BB: out_word = 8'h00;
		16'hB0BC: out_word = 8'hB7;
		16'hB0BD: out_word = 8'h28;
		16'hB0BE: out_word = 8'h04;
		16'hB0BF: out_word = 8'h19;
		16'hB0C0: out_word = 8'h3D;
		16'hB0C1: out_word = 8'h18;
		16'hB0C2: out_word = 8'hF9;
		16'hB0C3: out_word = 8'hEB;
		16'hB0C4: out_word = 8'hF1;
		16'hB0C5: out_word = 8'hC9;
		16'hB0C6: out_word = 8'hD5;
		16'hB0C7: out_word = 8'hCD;
		16'hB0C8: out_word = 8'hB4;
		16'hB0C9: out_word = 8'h30;
		16'hB0CA: out_word = 8'h26;
		16'hB0CB: out_word = 8'h00;
		16'hB0CC: out_word = 8'h68;
		16'hB0CD: out_word = 8'h19;
		16'hB0CE: out_word = 8'hD1;
		16'hB0CF: out_word = 8'hC9;
		16'hB0D0: out_word = 8'h05;
		16'hB0D1: out_word = 8'h00;
		16'hB0D2: out_word = 8'h00;
		16'hB0D3: out_word = 8'h00;
		16'hB0D4: out_word = 8'hF8;
		16'hB0D5: out_word = 8'hF6;
		16'hB0D6: out_word = 8'h21;
		16'hB0D7: out_word = 8'hD0;
		16'hB0D8: out_word = 8'h30;
		16'hB0D9: out_word = 8'h11;
		16'hB0DA: out_word = 8'hF5;
		16'hB0DB: out_word = 8'hF6;
		16'hB0DC: out_word = 8'hC3;
		16'hB0DD: out_word = 8'hBA;
		16'hB0DE: out_word = 8'h3F;
		16'hB0DF: out_word = 8'hC5;
		16'hB0E0: out_word = 8'hD5;
		16'hB0E1: out_word = 8'h21;
		16'hB0E2: out_word = 8'hF5;
		16'hB0E3: out_word = 8'hF6;
		16'hB0E4: out_word = 8'hE5;
		16'hB0E5: out_word = 8'h7E;
		16'hB0E6: out_word = 8'hB7;
		16'hB0E7: out_word = 8'h20;
		16'hB0E8: out_word = 8'h18;
		16'hB0E9: out_word = 8'hE5;
		16'hB0EA: out_word = 8'hCD;
		16'hB0EB: out_word = 8'h5F;
		16'hB0EC: out_word = 8'h33;
		16'hB0ED: out_word = 8'h2A;
		16'hB0EE: out_word = 8'hD7;
		16'hB0EF: out_word = 8'hF9;
		16'hB0F0: out_word = 8'hCD;
		16'hB0F1: out_word = 8'h52;
		16'hB0F2: out_word = 8'h33;
		16'hB0F3: out_word = 8'h30;
		16'hB0F4: out_word = 8'h03;
		16'hB0F5: out_word = 8'h22;
		16'hB0F6: out_word = 8'hD7;
		16'hB0F7: out_word = 8'hF9;
		16'hB0F8: out_word = 8'h44;
		16'hB0F9: out_word = 8'h4D;
		16'hB0FA: out_word = 8'hE1;
		16'hB0FB: out_word = 8'hCD;
		16'hB0FC: out_word = 8'hD6;
		16'hB0FD: out_word = 8'h32;
		16'hB0FE: out_word = 8'h3D;
		16'hB0FF: out_word = 8'h18;
		16'hB100: out_word = 8'h15;
		16'hB101: out_word = 8'h21;
		16'hB102: out_word = 8'h0D;
		16'hB103: out_word = 8'hEC;
		16'hB104: out_word = 8'hCB;
		16'hB105: out_word = 8'h86;
		16'hB106: out_word = 8'h21;
		16'hB107: out_word = 8'hF8;
		16'hB108: out_word = 8'hF6;
		16'hB109: out_word = 8'h54;
		16'hB10A: out_word = 8'h5D;
		16'hB10B: out_word = 8'h01;
		16'hB10C: out_word = 8'h23;
		16'hB10D: out_word = 8'h00;
		16'hB10E: out_word = 8'h09;
		16'hB10F: out_word = 8'h01;
		16'hB110: out_word = 8'hBC;
		16'hB111: out_word = 8'h02;
		16'hB112: out_word = 8'hED;
		16'hB113: out_word = 8'hB0;
		16'hB114: out_word = 8'h3D;
		16'hB115: out_word = 8'h37;
		16'hB116: out_word = 8'hD1;
		16'hB117: out_word = 8'h12;
		16'hB118: out_word = 8'h21;
		16'hB119: out_word = 8'hF8;
		16'hB11A: out_word = 8'hF6;
		16'hB11B: out_word = 8'hD1;
		16'hB11C: out_word = 8'hC1;
		16'hB11D: out_word = 8'hC9;
		16'hB11E: out_word = 8'hC5;
		16'hB11F: out_word = 8'hD5;
		16'hB120: out_word = 8'h21;
		16'hB121: out_word = 8'h20;
		16'hB122: out_word = 8'h00;
		16'hB123: out_word = 8'h19;
		16'hB124: out_word = 8'h7E;
		16'hB125: out_word = 8'h2F;
		16'hB126: out_word = 8'hE6;
		16'hB127: out_word = 8'h11;
		16'hB128: out_word = 8'h20;
		16'hB129: out_word = 8'h15;
		16'hB12A: out_word = 8'hE5;
		16'hB12B: out_word = 8'hD5;
		16'hB12C: out_word = 8'h23;
		16'hB12D: out_word = 8'h56;
		16'hB12E: out_word = 8'h23;
		16'hB12F: out_word = 8'h5E;
		16'hB130: out_word = 8'hD5;
		16'hB131: out_word = 8'hCD;
		16'hB132: out_word = 8'h5F;
		16'hB133: out_word = 8'h33;
		16'hB134: out_word = 8'hE1;
		16'hB135: out_word = 8'hCD;
		16'hB136: out_word = 8'h4A;
		16'hB137: out_word = 8'h33;
		16'hB138: out_word = 8'h30;
		16'hB139: out_word = 8'h03;
		16'hB13A: out_word = 8'h22;
		16'hB13B: out_word = 8'hD7;
		16'hB13C: out_word = 8'hF9;
		16'hB13D: out_word = 8'hD1;
		16'hB13E: out_word = 8'hE1;
		16'hB13F: out_word = 8'hCB;
		16'hB140: out_word = 8'h46;
		16'hB141: out_word = 8'h21;
		16'hB142: out_word = 8'hF5;
		16'hB143: out_word = 8'hF6;
		16'hB144: out_word = 8'hE5;
		16'hB145: out_word = 8'h28;
		16'hB146: out_word = 8'h05;
		16'hB147: out_word = 8'h3E;
		16'hB148: out_word = 8'h00;
		16'hB149: out_word = 8'h37;
		16'hB14A: out_word = 8'h18;
		16'hB14B: out_word = 8'hCA;
		16'hB14C: out_word = 8'h7E;
		16'hB14D: out_word = 8'hFE;
		16'hB14E: out_word = 8'h14;
		16'hB14F: out_word = 8'h28;
		16'hB150: out_word = 8'hC5;
		16'hB151: out_word = 8'h01;
		16'hB152: out_word = 8'h23;
		16'hB153: out_word = 8'h00;
		16'hB154: out_word = 8'h21;
		16'hB155: out_word = 8'hF8;
		16'hB156: out_word = 8'hF6;
		16'hB157: out_word = 8'hEB;
		16'hB158: out_word = 8'hED;
		16'hB159: out_word = 8'hB0;
		16'hB15A: out_word = 8'h21;
		16'hB15B: out_word = 8'hD6;
		16'hB15C: out_word = 8'hF9;
		16'hB15D: out_word = 8'h54;
		16'hB15E: out_word = 8'h5D;
		16'hB15F: out_word = 8'h01;
		16'hB160: out_word = 8'h23;
		16'hB161: out_word = 8'h00;
		16'hB162: out_word = 8'hB7;
		16'hB163: out_word = 8'hED;
		16'hB164: out_word = 8'h42;
		16'hB165: out_word = 8'h01;
		16'hB166: out_word = 8'hBC;
		16'hB167: out_word = 8'h02;
		16'hB168: out_word = 8'hED;
		16'hB169: out_word = 8'hB8;
		16'hB16A: out_word = 8'h3C;
		16'hB16B: out_word = 8'h37;
		16'hB16C: out_word = 8'h18;
		16'hB16D: out_word = 8'hA8;
		16'hB16E: out_word = 8'hC5;
		16'hB16F: out_word = 8'hD5;
		16'hB170: out_word = 8'hF5;
		16'hB171: out_word = 8'h06;
		16'hB172: out_word = 8'h00;
		16'hB173: out_word = 8'h0E;
		16'hB174: out_word = 8'h01;
		16'hB175: out_word = 8'hE5;
		16'hB176: out_word = 8'hCD;
		16'hB177: out_word = 8'hC3;
		16'hB178: out_word = 8'h31;
		16'hB179: out_word = 8'hE1;
		16'hB17A: out_word = 8'hCB;
		16'hB17B: out_word = 8'h5E;
		16'hB17C: out_word = 8'hCB;
		16'hB17D: out_word = 8'h9E;
		16'hB17E: out_word = 8'h20;
		16'hB17F: out_word = 8'h20;
		16'hB180: out_word = 8'hCD;
		16'hB181: out_word = 8'h41;
		16'hB182: out_word = 8'h2E;
		16'hB183: out_word = 8'hF1;
		16'hB184: out_word = 8'hCD;
		16'hB185: out_word = 8'hAC;
		16'hB186: out_word = 8'h16;
		16'hB187: out_word = 8'h28;
		16'hB188: out_word = 8'h31;
		16'hB189: out_word = 8'hF5;
		16'hB18A: out_word = 8'h06;
		16'hB18B: out_word = 8'h00;
		16'hB18C: out_word = 8'h0C;
		16'hB18D: out_word = 8'h79;
		16'hB18E: out_word = 8'hFE;
		16'hB18F: out_word = 8'h15;
		16'hB190: out_word = 8'h38;
		16'hB191: out_word = 8'h0E;
		16'hB192: out_word = 8'h2B;
		16'hB193: out_word = 8'h7E;
		16'hB194: out_word = 8'h23;
		16'hB195: out_word = 8'hFE;
		16'hB196: out_word = 8'h00;
		16'hB197: out_word = 8'h28;
		16'hB198: out_word = 8'h07;
		16'hB199: out_word = 8'hE5;
		16'hB19A: out_word = 8'h21;
		16'hB19B: out_word = 8'h0D;
		16'hB19C: out_word = 8'hEC;
		16'hB19D: out_word = 8'hCB;
		16'hB19E: out_word = 8'hC6;
		16'hB19F: out_word = 8'hE1;
		16'hB1A0: out_word = 8'hCB;
		16'hB1A1: out_word = 8'h4E;
		16'hB1A2: out_word = 8'hCB;
		16'hB1A3: out_word = 8'hCE;
		16'hB1A4: out_word = 8'hCB;
		16'hB1A5: out_word = 8'h9E;
		16'hB1A6: out_word = 8'hCD;
		16'hB1A7: out_word = 8'hC3;
		16'hB1A8: out_word = 8'h31;
		16'hB1A9: out_word = 8'h20;
		16'hB1AA: out_word = 8'hD5;
		16'hB1AB: out_word = 8'hC5;
		16'hB1AC: out_word = 8'hD5;
		16'hB1AD: out_word = 8'hCD;
		16'hB1AE: out_word = 8'hE6;
		16'hB1AF: out_word = 8'h35;
		16'hB1B0: out_word = 8'h36;
		16'hB1B1: out_word = 8'h08;
		16'hB1B2: out_word = 8'hD1;
		16'hB1B3: out_word = 8'hC1;
		16'hB1B4: out_word = 8'hCD;
		16'hB1B5: out_word = 8'hF4;
		16'hB1B6: out_word = 8'h35;
		16'hB1B7: out_word = 8'hF1;
		16'hB1B8: out_word = 8'h18;
		16'hB1B9: out_word = 8'hCA;
		16'hB1BA: out_word = 8'h79;
		16'hB1BB: out_word = 8'h32;
		16'hB1BC: out_word = 8'hF5;
		16'hB1BD: out_word = 8'hF6;
		16'hB1BE: out_word = 8'hCB;
		16'hB1BF: out_word = 8'hDE;
		16'hB1C0: out_word = 8'hD1;
		16'hB1C1: out_word = 8'hC1;
		16'hB1C2: out_word = 8'hC9;
		16'hB1C3: out_word = 8'h21;
		16'hB1C4: out_word = 8'hF8;
		16'hB1C5: out_word = 8'hF6;
		16'hB1C6: out_word = 8'hC3;
		16'hB1C7: out_word = 8'hB7;
		16'hB1C8: out_word = 8'h30;
		16'hB1C9: out_word = 8'hC5;
		16'hB1CA: out_word = 8'hD5;
		16'hB1CB: out_word = 8'h21;
		16'hB1CC: out_word = 8'h0D;
		16'hB1CD: out_word = 8'hEC;
		16'hB1CE: out_word = 8'hCB;
		16'hB1CF: out_word = 8'h86;
		16'hB1D0: out_word = 8'h3A;
		16'hB1D1: out_word = 8'hF5;
		16'hB1D2: out_word = 8'hF6;
		16'hB1D3: out_word = 8'h4F;
		16'hB1D4: out_word = 8'hB7;
		16'hB1D5: out_word = 8'h3E;
		16'hB1D6: out_word = 8'h00;
		16'hB1D7: out_word = 8'h28;
		16'hB1D8: out_word = 8'h42;
		16'hB1D9: out_word = 8'hCD;
		16'hB1DA: out_word = 8'hC3;
		16'hB1DB: out_word = 8'h31;
		16'hB1DC: out_word = 8'hF5;
		16'hB1DD: out_word = 8'h06;
		16'hB1DE: out_word = 8'h00;
		16'hB1DF: out_word = 8'hCD;
		16'hB1E0: out_word = 8'h41;
		16'hB1E1: out_word = 8'h2E;
		16'hB1E2: out_word = 8'h30;
		16'hB1E3: out_word = 8'h0E;
		16'hB1E4: out_word = 8'hF1;
		16'hB1E5: out_word = 8'hCD;
		16'hB1E6: out_word = 8'hC1;
		16'hB1E7: out_word = 8'h16;
		16'hB1E8: out_word = 8'hF5;
		16'hB1E9: out_word = 8'hC5;
		16'hB1EA: out_word = 8'h06;
		16'hB1EB: out_word = 8'h00;
		16'hB1EC: out_word = 8'hCD;
		16'hB1ED: out_word = 8'h41;
		16'hB1EE: out_word = 8'h2E;
		16'hB1EF: out_word = 8'hC1;
		16'hB1F0: out_word = 8'h38;
		16'hB1F1: out_word = 8'h24;
		16'hB1F2: out_word = 8'h23;
		16'hB1F3: out_word = 8'h7E;
		16'hB1F4: out_word = 8'hF5;
		16'hB1F5: out_word = 8'hC5;
		16'hB1F6: out_word = 8'h79;
		16'hB1F7: out_word = 8'hFE;
		16'hB1F8: out_word = 8'h01;
		16'hB1F9: out_word = 8'h20;
		16'hB1FA: out_word = 8'h09;
		16'hB1FB: out_word = 8'h3A;
		16'hB1FC: out_word = 8'h15;
		16'hB1FD: out_word = 8'hEC;
		16'hB1FE: out_word = 8'h4F;
		16'hB1FF: out_word = 8'hCD;
		16'hB200: out_word = 8'hB4;
		16'hB201: out_word = 8'h30;
		16'hB202: out_word = 8'h18;
		16'hB203: out_word = 8'h04;
		16'hB204: out_word = 8'h0D;
		16'hB205: out_word = 8'hCD;
		16'hB206: out_word = 8'hC3;
		16'hB207: out_word = 8'h31;
		16'hB208: out_word = 8'hC1;
		16'hB209: out_word = 8'hF1;
		16'hB20A: out_word = 8'h21;
		16'hB20B: out_word = 8'h20;
		16'hB20C: out_word = 8'h00;
		16'hB20D: out_word = 8'h19;
		16'hB20E: out_word = 8'hCB;
		16'hB20F: out_word = 8'h8E;
		16'hB210: out_word = 8'hB6;
		16'hB211: out_word = 8'h77;
		16'hB212: out_word = 8'h21;
		16'hB213: out_word = 8'hF5;
		16'hB214: out_word = 8'hF6;
		16'hB215: out_word = 8'h35;
		16'hB216: out_word = 8'hF1;
		16'hB217: out_word = 8'h0D;
		16'hB218: out_word = 8'h20;
		16'hB219: out_word = 8'hBF;
		16'hB21A: out_word = 8'h37;
		16'hB21B: out_word = 8'hD1;
		16'hB21C: out_word = 8'hC1;
		16'hB21D: out_word = 8'hC9;
		16'hB21E: out_word = 8'h03;
		16'hB21F: out_word = 8'h00;
		16'hB220: out_word = 8'hDE;
		16'hB221: out_word = 8'hF9;
		16'hB222: out_word = 8'h21;
		16'hB223: out_word = 8'h1E;
		16'hB224: out_word = 8'h32;
		16'hB225: out_word = 8'h11;
		16'hB226: out_word = 8'hDB;
		16'hB227: out_word = 8'hF9;
		16'hB228: out_word = 8'hC3;
		16'hB229: out_word = 8'hBA;
		16'hB22A: out_word = 8'h3F;
		16'hB22B: out_word = 8'hC5;
		16'hB22C: out_word = 8'hD5;
		16'hB22D: out_word = 8'h21;
		16'hB22E: out_word = 8'hDB;
		16'hB22F: out_word = 8'hF9;
		16'hB230: out_word = 8'hE5;
		16'hB231: out_word = 8'h7E;
		16'hB232: out_word = 8'hB7;
		16'hB233: out_word = 8'h20;
		16'hB234: out_word = 8'h1E;
		16'hB235: out_word = 8'hE5;
		16'hB236: out_word = 8'hCD;
		16'hB237: out_word = 8'h5F;
		16'hB238: out_word = 8'h33;
		16'hB239: out_word = 8'h2A;
		16'hB23A: out_word = 8'h9A;
		16'hB23B: out_word = 8'hFC;
		16'hB23C: out_word = 8'hCD;
		16'hB23D: out_word = 8'h4A;
		16'hB23E: out_word = 8'h33;
		16'hB23F: out_word = 8'h30;
		16'hB240: out_word = 8'h03;
		16'hB241: out_word = 8'h22;
		16'hB242: out_word = 8'h9A;
		16'hB243: out_word = 8'hFC;
		16'hB244: out_word = 8'h44;
		16'hB245: out_word = 8'h4D;
		16'hB246: out_word = 8'hE1;
		16'hB247: out_word = 8'h23;
		16'hB248: out_word = 8'h23;
		16'hB249: out_word = 8'h23;
		16'hB24A: out_word = 8'h30;
		16'hB24B: out_word = 8'h11;
		16'hB24C: out_word = 8'hCD;
		16'hB24D: out_word = 8'hD6;
		16'hB24E: out_word = 8'h32;
		16'hB24F: out_word = 8'h3D;
		16'hB250: out_word = 8'hEB;
		16'hB251: out_word = 8'h18;
		16'hB252: out_word = 8'h0A;
		16'hB253: out_word = 8'h2A;
		16'hB254: out_word = 8'hDC;
		16'hB255: out_word = 8'hF9;
		16'hB256: out_word = 8'h01;
		16'hB257: out_word = 8'h23;
		16'hB258: out_word = 8'h00;
		16'hB259: out_word = 8'hED;
		16'hB25A: out_word = 8'h42;
		16'hB25B: out_word = 8'h37;
		16'hB25C: out_word = 8'h3D;
		16'hB25D: out_word = 8'hEB;
		16'hB25E: out_word = 8'hE1;
		16'hB25F: out_word = 8'h30;
		16'hB260: out_word = 8'h01;
		16'hB261: out_word = 8'h77;
		16'hB262: out_word = 8'h23;
		16'hB263: out_word = 8'h73;
		16'hB264: out_word = 8'h23;
		16'hB265: out_word = 8'h72;
		16'hB266: out_word = 8'hEB;
		16'hB267: out_word = 8'hD1;
		16'hB268: out_word = 8'hC1;
		16'hB269: out_word = 8'hC9;
		16'hB26A: out_word = 8'hC5;
		16'hB26B: out_word = 8'hD5;
		16'hB26C: out_word = 8'h21;
		16'hB26D: out_word = 8'h20;
		16'hB26E: out_word = 8'h00;
		16'hB26F: out_word = 8'h19;
		16'hB270: out_word = 8'h7E;
		16'hB271: out_word = 8'h2F;
		16'hB272: out_word = 8'hE6;
		16'hB273: out_word = 8'h11;
		16'hB274: out_word = 8'h20;
		16'hB275: out_word = 8'h0C;
		16'hB276: out_word = 8'hD5;
		16'hB277: out_word = 8'hE5;
		16'hB278: out_word = 8'h23;
		16'hB279: out_word = 8'h56;
		16'hB27A: out_word = 8'h23;
		16'hB27B: out_word = 8'h5E;
		16'hB27C: out_word = 8'hED;
		16'hB27D: out_word = 8'h53;
		16'hB27E: out_word = 8'h9A;
		16'hB27F: out_word = 8'hFC;
		16'hB280: out_word = 8'hE1;
		16'hB281: out_word = 8'hD1;
		16'hB282: out_word = 8'hCB;
		16'hB283: out_word = 8'h5E;
		16'hB284: out_word = 8'h21;
		16'hB285: out_word = 8'hDB;
		16'hB286: out_word = 8'hF9;
		16'hB287: out_word = 8'hE5;
		16'hB288: out_word = 8'h28;
		16'hB289: out_word = 8'h16;
		16'hB28A: out_word = 8'hE5;
		16'hB28B: out_word = 8'hCD;
		16'hB28C: out_word = 8'h5F;
		16'hB28D: out_word = 8'h33;
		16'hB28E: out_word = 8'h2A;
		16'hB28F: out_word = 8'h9A;
		16'hB290: out_word = 8'hFC;
		16'hB291: out_word = 8'hCD;
		16'hB292: out_word = 8'h52;
		16'hB293: out_word = 8'h33;
		16'hB294: out_word = 8'h22;
		16'hB295: out_word = 8'h9A;
		16'hB296: out_word = 8'hFC;
		16'hB297: out_word = 8'hE1;
		16'hB298: out_word = 8'h23;
		16'hB299: out_word = 8'h23;
		16'hB29A: out_word = 8'h23;
		16'hB29B: out_word = 8'h3E;
		16'hB29C: out_word = 8'h00;
		16'hB29D: out_word = 8'h37;
		16'hB29E: out_word = 8'h18;
		16'hB29F: out_word = 8'hBD;
		16'hB2A0: out_word = 8'h7E;
		16'hB2A1: out_word = 8'hFE;
		16'hB2A2: out_word = 8'h14;
		16'hB2A3: out_word = 8'h28;
		16'hB2A4: out_word = 8'h0E;
		16'hB2A5: out_word = 8'h3C;
		16'hB2A6: out_word = 8'h2A;
		16'hB2A7: out_word = 8'hDC;
		16'hB2A8: out_word = 8'hF9;
		16'hB2A9: out_word = 8'h01;
		16'hB2AA: out_word = 8'h23;
		16'hB2AB: out_word = 8'h00;
		16'hB2AC: out_word = 8'hEB;
		16'hB2AD: out_word = 8'hED;
		16'hB2AE: out_word = 8'hB0;
		16'hB2AF: out_word = 8'hEB;
		16'hB2B0: out_word = 8'h37;
		16'hB2B1: out_word = 8'h18;
		16'hB2B2: out_word = 8'hAA;
		16'hB2B3: out_word = 8'hE1;
		16'hB2B4: out_word = 8'hD1;
		16'hB2B5: out_word = 8'hC1;
		16'hB2B6: out_word = 8'hC9;
		16'hB2B7: out_word = 8'h21;
		16'hB2B8: out_word = 8'hDE;
		16'hB2B9: out_word = 8'hF9;
		16'hB2BA: out_word = 8'hC3;
		16'hB2BB: out_word = 8'hB7;
		16'hB2BC: out_word = 8'h30;
		16'hB2BD: out_word = 8'h08;
		16'hB2BE: out_word = 8'h0D;
		16'hB2BF: out_word = 8'hCC;
		16'hB2C0: out_word = 8'h35;
		16'hB2C1: out_word = 8'h01;
		16'hB2C2: out_word = 8'hDA;
		16'hB2C3: out_word = 8'h35;
		16'hB2C4: out_word = 8'h12;
		16'hB2C5: out_word = 8'h5A;
		16'hB2C6: out_word = 8'h33;
		16'hB2C7: out_word = 8'h13;
		16'hB2C8: out_word = 8'h5A;
		16'hB2C9: out_word = 8'h33;
		16'hB2CA: out_word = 8'h14;
		16'hB2CB: out_word = 8'h5A;
		16'hB2CC: out_word = 8'h33;
		16'hB2CD: out_word = 8'h15;
		16'hB2CE: out_word = 8'h5A;
		16'hB2CF: out_word = 8'h33;
		16'hB2D0: out_word = 8'h10;
		16'hB2D1: out_word = 8'h5A;
		16'hB2D2: out_word = 8'h33;
		16'hB2D3: out_word = 8'h11;
		16'hB2D4: out_word = 8'h5A;
		16'hB2D5: out_word = 8'h33;
		16'hB2D6: out_word = 8'h54;
		16'hB2D7: out_word = 8'h5D;
		16'hB2D8: out_word = 8'h13;
		16'hB2D9: out_word = 8'h13;
		16'hB2DA: out_word = 8'h13;
		16'hB2DB: out_word = 8'hD5;
		16'hB2DC: out_word = 8'h21;
		16'hB2DD: out_word = 8'h20;
		16'hB2DE: out_word = 8'h00;
		16'hB2DF: out_word = 8'h19;
		16'hB2E0: out_word = 8'h36;
		16'hB2E1: out_word = 8'h01;
		16'hB2E2: out_word = 8'h23;
		16'hB2E3: out_word = 8'h70;
		16'hB2E4: out_word = 8'h23;
		16'hB2E5: out_word = 8'h71;
		16'hB2E6: out_word = 8'h0E;
		16'hB2E7: out_word = 8'h01;
		16'hB2E8: out_word = 8'h06;
		16'hB2E9: out_word = 8'h00;
		16'hB2EA: out_word = 8'hC5;
		16'hB2EB: out_word = 8'hD5;
		16'hB2EC: out_word = 8'h3A;
		16'hB2ED: out_word = 8'h0E;
		16'hB2EE: out_word = 8'hEC;
		16'hB2EF: out_word = 8'hFE;
		16'hB2F0: out_word = 8'h04;
		16'hB2F1: out_word = 8'hC4;
		16'hB2F2: out_word = 8'h17;
		16'hB2F3: out_word = 8'h35;
		16'hB2F4: out_word = 8'hD1;
		16'hB2F5: out_word = 8'hC1;
		16'hB2F6: out_word = 8'h38;
		16'hB2F7: out_word = 8'h0F;
		16'hB2F8: out_word = 8'h79;
		16'hB2F9: out_word = 8'hFE;
		16'hB2FA: out_word = 8'h01;
		16'hB2FB: out_word = 8'h3E;
		16'hB2FC: out_word = 8'h0D;
		16'hB2FD: out_word = 8'h20;
		16'hB2FE: out_word = 8'h08;
		16'hB2FF: out_word = 8'h78;
		16'hB300: out_word = 8'hB7;
		16'hB301: out_word = 8'h3E;
		16'hB302: out_word = 8'h01;
		16'hB303: out_word = 8'h28;
		16'hB304: out_word = 8'h02;
		16'hB305: out_word = 8'h3E;
		16'hB306: out_word = 8'h0D;
		16'hB307: out_word = 8'h21;
		16'hB308: out_word = 8'hBD;
		16'hB309: out_word = 8'h32;
		16'hB30A: out_word = 8'hCD;
		16'hB30B: out_word = 8'hCE;
		16'hB30C: out_word = 8'h3F;
		16'hB30D: out_word = 8'h38;
		16'hB30E: out_word = 8'h1D;
		16'hB30F: out_word = 8'h28;
		16'hB310: out_word = 8'hD9;
		16'hB311: out_word = 8'hF5;
		16'hB312: out_word = 8'h3E;
		16'hB313: out_word = 8'h1F;
		16'hB314: out_word = 8'hB8;
		16'hB315: out_word = 8'h30;
		16'hB316: out_word = 8'h0F;
		16'hB317: out_word = 8'h3E;
		16'hB318: out_word = 8'h12;
		16'hB319: out_word = 8'hCD;
		16'hB31A: out_word = 8'h31;
		16'hB31B: out_word = 8'h33;
		16'hB31C: out_word = 8'h38;
		16'hB31D: out_word = 8'h05;
		16'hB31E: out_word = 8'hF1;
		16'hB31F: out_word = 8'h3E;
		16'hB320: out_word = 8'h0D;
		16'hB321: out_word = 8'h18;
		16'hB322: out_word = 8'hE4;
		16'hB323: out_word = 8'hCD;
		16'hB324: out_word = 8'hF4;
		16'hB325: out_word = 8'h35;
		16'hB326: out_word = 8'hF1;
		16'hB327: out_word = 8'hCD;
		16'hB328: out_word = 8'hC5;
		16'hB329: out_word = 8'h35;
		16'hB32A: out_word = 8'h18;
		16'hB32B: out_word = 8'hBE;
		16'hB32C: out_word = 8'hE1;
		16'hB32D: out_word = 8'h79;
		16'hB32E: out_word = 8'hC8;
		16'hB32F: out_word = 8'h37;
		16'hB330: out_word = 8'hC9;
		16'hB331: out_word = 8'hF5;
		16'hB332: out_word = 8'hCD;
		16'hB333: out_word = 8'hE6;
		16'hB334: out_word = 8'h35;
		16'hB335: out_word = 8'hF1;
		16'hB336: out_word = 8'hAE;
		16'hB337: out_word = 8'h77;
		16'hB338: out_word = 8'h79;
		16'hB339: out_word = 8'hFE;
		16'hB33A: out_word = 8'h14;
		16'hB33B: out_word = 8'hD0;
		16'hB33C: out_word = 8'h0C;
		16'hB33D: out_word = 8'h21;
		16'hB33E: out_word = 8'h23;
		16'hB33F: out_word = 8'h00;
		16'hB340: out_word = 8'h19;
		16'hB341: out_word = 8'hEB;
		16'hB342: out_word = 8'h21;
		16'hB343: out_word = 8'h20;
		16'hB344: out_word = 8'h00;
		16'hB345: out_word = 8'h19;
		16'hB346: out_word = 8'h36;
		16'hB347: out_word = 8'h00;
		16'hB348: out_word = 8'h37;
		16'hB349: out_word = 8'hC9;
		16'hB34A: out_word = 8'hCD;
		16'hB34B: out_word = 8'hB6;
		16'hB34C: out_word = 8'h34;
		16'hB34D: out_word = 8'hD8;
		16'hB34E: out_word = 8'h21;
		16'hB34F: out_word = 8'h00;
		16'hB350: out_word = 8'h00;
		16'hB351: out_word = 8'hC9;
		16'hB352: out_word = 8'hCD;
		16'hB353: out_word = 8'h30;
		16'hB354: out_word = 8'h34;
		16'hB355: out_word = 8'hD8;
		16'hB356: out_word = 8'h21;
		16'hB357: out_word = 8'h00;
		16'hB358: out_word = 8'h00;
		16'hB359: out_word = 8'hC9;
		16'hB35A: out_word = 8'hCD;
		16'hB35B: out_word = 8'h17;
		16'hB35C: out_word = 8'h35;
		16'hB35D: out_word = 8'h3F;
		16'hB35E: out_word = 8'hD0;
		16'hB35F: out_word = 8'h21;
		16'hB360: out_word = 8'h00;
		16'hB361: out_word = 8'h00;
		16'hB362: out_word = 8'h22;
		16'hB363: out_word = 8'h9F;
		16'hB364: out_word = 8'hFC;
		16'hB365: out_word = 8'h22;
		16'hB366: out_word = 8'hA1;
		16'hB367: out_word = 8'hFC;
		16'hB368: out_word = 8'h21;
		16'hB369: out_word = 8'h74;
		16'hB36A: out_word = 8'h33;
		16'hB36B: out_word = 8'h11;
		16'hB36C: out_word = 8'hAE;
		16'hB36D: out_word = 8'hFC;
		16'hB36E: out_word = 8'h01;
		16'hB36F: out_word = 8'hBC;
		16'hB370: out_word = 8'h00;
		16'hB371: out_word = 8'hED;
		16'hB372: out_word = 8'hB0;
		16'hB373: out_word = 8'hC9;
		16'hB374: out_word = 8'hF3;
		16'hB375: out_word = 8'h01;
		16'hB376: out_word = 8'hFD;
		16'hB377: out_word = 8'h7F;
		16'hB378: out_word = 8'h16;
		16'hB379: out_word = 8'h17;
		16'hB37A: out_word = 8'hED;
		16'hB37B: out_word = 8'h51;
		16'hB37C: out_word = 8'hFE;
		16'hB37D: out_word = 8'h50;
		16'hB37E: out_word = 8'h30;
		16'hB37F: out_word = 8'h31;
		16'hB380: out_word = 8'hFE;
		16'hB381: out_word = 8'h40;
		16'hB382: out_word = 8'h30;
		16'hB383: out_word = 8'h26;
		16'hB384: out_word = 8'hFE;
		16'hB385: out_word = 8'h30;
		16'hB386: out_word = 8'h30;
		16'hB387: out_word = 8'h1B;
		16'hB388: out_word = 8'hFE;
		16'hB389: out_word = 8'h20;
		16'hB38A: out_word = 8'h30;
		16'hB38B: out_word = 8'h10;
		16'hB38C: out_word = 8'hFE;
		16'hB38D: out_word = 8'h10;
		16'hB38E: out_word = 8'h30;
		16'hB38F: out_word = 8'h05;
		16'hB390: out_word = 8'h21;
		16'hB391: out_word = 8'h96;
		16'hB392: out_word = 8'h00;
		16'hB393: out_word = 8'h18;
		16'hB394: out_word = 8'h21;
		16'hB395: out_word = 8'hD6;
		16'hB396: out_word = 8'h10;
		16'hB397: out_word = 8'h21;
		16'hB398: out_word = 8'hCF;
		16'hB399: out_word = 8'h00;
		16'hB39A: out_word = 8'h18;
		16'hB39B: out_word = 8'h1A;
		16'hB39C: out_word = 8'hD6;
		16'hB39D: out_word = 8'h20;
		16'hB39E: out_word = 8'h21;
		16'hB39F: out_word = 8'h00;
		16'hB3A0: out_word = 8'h01;
		16'hB3A1: out_word = 8'h18;
		16'hB3A2: out_word = 8'h13;
		16'hB3A3: out_word = 8'hD6;
		16'hB3A4: out_word = 8'h30;
		16'hB3A5: out_word = 8'h21;
		16'hB3A6: out_word = 8'h3E;
		16'hB3A7: out_word = 8'h01;
		16'hB3A8: out_word = 8'h18;
		16'hB3A9: out_word = 8'h0C;
		16'hB3AA: out_word = 8'hD6;
		16'hB3AB: out_word = 8'h40;
		16'hB3AC: out_word = 8'h21;
		16'hB3AD: out_word = 8'h8B;
		16'hB3AE: out_word = 8'h01;
		16'hB3AF: out_word = 8'h18;
		16'hB3B0: out_word = 8'h05;
		16'hB3B1: out_word = 8'hD6;
		16'hB3B2: out_word = 8'h50;
		16'hB3B3: out_word = 8'h21;
		16'hB3B4: out_word = 8'hD4;
		16'hB3B5: out_word = 8'h01;
		16'hB3B6: out_word = 8'h47;
		16'hB3B7: out_word = 8'hB7;
		16'hB3B8: out_word = 8'h28;
		16'hB3B9: out_word = 8'h09;
		16'hB3BA: out_word = 8'h7E;
		16'hB3BB: out_word = 8'h23;
		16'hB3BC: out_word = 8'hE6;
		16'hB3BD: out_word = 8'h80;
		16'hB3BE: out_word = 8'h28;
		16'hB3BF: out_word = 8'hFA;
		16'hB3C0: out_word = 8'h05;
		16'hB3C1: out_word = 8'h18;
		16'hB3C2: out_word = 8'hF5;
		16'hB3C3: out_word = 8'h11;
		16'hB3C4: out_word = 8'hA3;
		16'hB3C5: out_word = 8'hFC;
		16'hB3C6: out_word = 8'hED;
		16'hB3C7: out_word = 8'h53;
		16'hB3C8: out_word = 8'hA1;
		16'hB3C9: out_word = 8'hFC;
		16'hB3CA: out_word = 8'h3A;
		16'hB3CB: out_word = 8'h9E;
		16'hB3CC: out_word = 8'hFC;
		16'hB3CD: out_word = 8'hB7;
		16'hB3CE: out_word = 8'h3E;
		16'hB3CF: out_word = 8'h00;
		16'hB3D0: out_word = 8'h32;
		16'hB3D1: out_word = 8'h9E;
		16'hB3D2: out_word = 8'hFC;
		16'hB3D3: out_word = 8'h20;
		16'hB3D4: out_word = 8'h04;
		16'hB3D5: out_word = 8'h3E;
		16'hB3D6: out_word = 8'h20;
		16'hB3D7: out_word = 8'h12;
		16'hB3D8: out_word = 8'h13;
		16'hB3D9: out_word = 8'h7E;
		16'hB3DA: out_word = 8'h47;
		16'hB3DB: out_word = 8'h23;
		16'hB3DC: out_word = 8'h12;
		16'hB3DD: out_word = 8'h13;
		16'hB3DE: out_word = 8'hE6;
		16'hB3DF: out_word = 8'h80;
		16'hB3E0: out_word = 8'h28;
		16'hB3E1: out_word = 8'hF7;
		16'hB3E2: out_word = 8'h78;
		16'hB3E3: out_word = 8'hE6;
		16'hB3E4: out_word = 8'h7F;
		16'hB3E5: out_word = 8'h1B;
		16'hB3E6: out_word = 8'h12;
		16'hB3E7: out_word = 8'h13;
		16'hB3E8: out_word = 8'h3E;
		16'hB3E9: out_word = 8'hA0;
		16'hB3EA: out_word = 8'h12;
		16'hB3EB: out_word = 8'h3E;
		16'hB3EC: out_word = 8'h07;
		16'hB3ED: out_word = 8'h01;
		16'hB3EE: out_word = 8'hFD;
		16'hB3EF: out_word = 8'h7F;
		16'hB3F0: out_word = 8'hED;
		16'hB3F1: out_word = 8'h79;
		16'hB3F2: out_word = 8'hFB;
		16'hB3F3: out_word = 8'hC9;
		16'hB3F4: out_word = 8'hF3;
		16'hB3F5: out_word = 8'h01;
		16'hB3F6: out_word = 8'hFD;
		16'hB3F7: out_word = 8'h7F;
		16'hB3F8: out_word = 8'h16;
		16'hB3F9: out_word = 8'h17;
		16'hB3FA: out_word = 8'hED;
		16'hB3FB: out_word = 8'h51;
		16'hB3FC: out_word = 8'h21;
		16'hB3FD: out_word = 8'h96;
		16'hB3FE: out_word = 8'h00;
		16'hB3FF: out_word = 8'h06;
		16'hB400: out_word = 8'hA5;
		16'hB401: out_word = 8'h11;
		16'hB402: out_word = 8'h74;
		16'hB403: out_word = 8'hFD;
		16'hB404: out_word = 8'h1A;
		16'hB405: out_word = 8'hE6;
		16'hB406: out_word = 8'h7F;
		16'hB407: out_word = 8'hFE;
		16'hB408: out_word = 8'h61;
		16'hB409: out_word = 8'h1A;
		16'hB40A: out_word = 8'h38;
		16'hB40B: out_word = 8'h02;
		16'hB40C: out_word = 8'hE6;
		16'hB40D: out_word = 8'hDF;
		16'hB40E: out_word = 8'hBE;
		16'hB40F: out_word = 8'h20;
		16'hB410: out_word = 8'h09;
		16'hB411: out_word = 8'h23;
		16'hB412: out_word = 8'h13;
		16'hB413: out_word = 8'hE6;
		16'hB414: out_word = 8'h80;
		16'hB415: out_word = 8'h28;
		16'hB416: out_word = 8'hED;
		16'hB417: out_word = 8'h37;
		16'hB418: out_word = 8'h18;
		16'hB419: out_word = 8'h0C;
		16'hB41A: out_word = 8'h04;
		16'hB41B: out_word = 8'h28;
		16'hB41C: out_word = 8'h08;
		16'hB41D: out_word = 8'h7E;
		16'hB41E: out_word = 8'hE6;
		16'hB41F: out_word = 8'h80;
		16'hB420: out_word = 8'h23;
		16'hB421: out_word = 8'h28;
		16'hB422: out_word = 8'hFA;
		16'hB423: out_word = 8'h18;
		16'hB424: out_word = 8'hDC;
		16'hB425: out_word = 8'hB7;
		16'hB426: out_word = 8'h78;
		16'hB427: out_word = 8'h16;
		16'hB428: out_word = 8'h07;
		16'hB429: out_word = 8'h01;
		16'hB42A: out_word = 8'hFD;
		16'hB42B: out_word = 8'h7F;
		16'hB42C: out_word = 8'hED;
		16'hB42D: out_word = 8'h51;
		16'hB42E: out_word = 8'hFB;
		16'hB42F: out_word = 8'hC9;
		16'hB430: out_word = 8'hCD;
		16'hB431: out_word = 8'hEA;
		16'hB432: out_word = 8'h34;
		16'hB433: out_word = 8'hB7;
		16'hB434: out_word = 8'h32;
		16'hB435: out_word = 8'h9E;
		16'hB436: out_word = 8'hFC;
		16'hB437: out_word = 8'hCD;
		16'hB438: out_word = 8'h20;
		16'hB439: out_word = 8'h1F;
		16'hB43A: out_word = 8'hCD;
		16'hB43B: out_word = 8'hF6;
		16'hB43C: out_word = 8'h34;
		16'hB43D: out_word = 8'h30;
		16'hB43E: out_word = 8'h52;
		16'hB43F: out_word = 8'h20;
		16'hB440: out_word = 8'h0C;
		16'hB441: out_word = 8'h78;
		16'hB442: out_word = 8'hB1;
		16'hB443: out_word = 8'h28;
		16'hB444: out_word = 8'h08;
		16'hB445: out_word = 8'hCD;
		16'hB446: out_word = 8'hCF;
		16'hB447: out_word = 8'h34;
		16'hB448: out_word = 8'hCD;
		16'hB449: out_word = 8'hD9;
		16'hB44A: out_word = 8'h34;
		16'hB44B: out_word = 8'h30;
		16'hB44C: out_word = 8'h44;
		16'hB44D: out_word = 8'h56;
		16'hB44E: out_word = 8'h23;
		16'hB44F: out_word = 8'h5E;
		16'hB450: out_word = 8'hCD;
		16'hB451: out_word = 8'h45;
		16'hB452: out_word = 8'h1F;
		16'hB453: out_word = 8'hD5;
		16'hB454: out_word = 8'hE5;
		16'hB455: out_word = 8'hDD;
		16'hB456: out_word = 8'hE5;
		16'hB457: out_word = 8'hDD;
		16'hB458: out_word = 8'h21;
		16'hB459: out_word = 8'hA3;
		16'hB45A: out_word = 8'hFC;
		16'hB45B: out_word = 8'hDD;
		16'hB45C: out_word = 8'h22;
		16'hB45D: out_word = 8'hA1;
		16'hB45E: out_word = 8'hFC;
		16'hB45F: out_word = 8'hEB;
		16'hB460: out_word = 8'h06;
		16'hB461: out_word = 8'h00;
		16'hB462: out_word = 8'h11;
		16'hB463: out_word = 8'h18;
		16'hB464: out_word = 8'hFC;
		16'hB465: out_word = 8'hCD;
		16'hB466: out_word = 8'h95;
		16'hB467: out_word = 8'h34;
		16'hB468: out_word = 8'h11;
		16'hB469: out_word = 8'h9C;
		16'hB46A: out_word = 8'hFF;
		16'hB46B: out_word = 8'hCD;
		16'hB46C: out_word = 8'h95;
		16'hB46D: out_word = 8'h34;
		16'hB46E: out_word = 8'h11;
		16'hB46F: out_word = 8'hF6;
		16'hB470: out_word = 8'hFF;
		16'hB471: out_word = 8'hCD;
		16'hB472: out_word = 8'h95;
		16'hB473: out_word = 8'h34;
		16'hB474: out_word = 8'h11;
		16'hB475: out_word = 8'hFF;
		16'hB476: out_word = 8'hFF;
		16'hB477: out_word = 8'hCD;
		16'hB478: out_word = 8'h95;
		16'hB479: out_word = 8'h34;
		16'hB47A: out_word = 8'hDD;
		16'hB47B: out_word = 8'h2B;
		16'hB47C: out_word = 8'hDD;
		16'hB47D: out_word = 8'h7E;
		16'hB47E: out_word = 8'h00;
		16'hB47F: out_word = 8'hF6;
		16'hB480: out_word = 8'h80;
		16'hB481: out_word = 8'hDD;
		16'hB482: out_word = 8'h77;
		16'hB483: out_word = 8'h00;
		16'hB484: out_word = 8'hDD;
		16'hB485: out_word = 8'hE1;
		16'hB486: out_word = 8'hE1;
		16'hB487: out_word = 8'hD1;
		16'hB488: out_word = 8'h23;
		16'hB489: out_word = 8'h23;
		16'hB48A: out_word = 8'h23;
		16'hB48B: out_word = 8'h22;
		16'hB48C: out_word = 8'h9F;
		16'hB48D: out_word = 8'hFC;
		16'hB48E: out_word = 8'hEB;
		16'hB48F: out_word = 8'h37;
		16'hB490: out_word = 8'hC9;
		16'hB491: out_word = 8'hCD;
		16'hB492: out_word = 8'h45;
		16'hB493: out_word = 8'h1F;
		16'hB494: out_word = 8'hC9;
		16'hB495: out_word = 8'hAF;
		16'hB496: out_word = 8'h19;
		16'hB497: out_word = 8'h3C;
		16'hB498: out_word = 8'h38;
		16'hB499: out_word = 8'hFC;
		16'hB49A: out_word = 8'hED;
		16'hB49B: out_word = 8'h52;
		16'hB49C: out_word = 8'h3D;
		16'hB49D: out_word = 8'hC6;
		16'hB49E: out_word = 8'h30;
		16'hB49F: out_word = 8'hDD;
		16'hB4A0: out_word = 8'h77;
		16'hB4A1: out_word = 8'h00;
		16'hB4A2: out_word = 8'hFE;
		16'hB4A3: out_word = 8'h30;
		16'hB4A4: out_word = 8'h20;
		16'hB4A5: out_word = 8'h0B;
		16'hB4A6: out_word = 8'h78;
		16'hB4A7: out_word = 8'hB7;
		16'hB4A8: out_word = 8'h20;
		16'hB4A9: out_word = 8'h09;
		16'hB4AA: out_word = 8'h3E;
		16'hB4AB: out_word = 8'h00;
		16'hB4AC: out_word = 8'hDD;
		16'hB4AD: out_word = 8'h77;
		16'hB4AE: out_word = 8'h00;
		16'hB4AF: out_word = 8'h18;
		16'hB4B0: out_word = 8'h02;
		16'hB4B1: out_word = 8'h06;
		16'hB4B2: out_word = 8'h01;
		16'hB4B3: out_word = 8'hDD;
		16'hB4B4: out_word = 8'h23;
		16'hB4B5: out_word = 8'hC9;
		16'hB4B6: out_word = 8'hCD;
		16'hB4B7: out_word = 8'hEA;
		16'hB4B8: out_word = 8'h34;
		16'hB4B9: out_word = 8'hB7;
		16'hB4BA: out_word = 8'h32;
		16'hB4BB: out_word = 8'h9E;
		16'hB4BC: out_word = 8'hFC;
		16'hB4BD: out_word = 8'hCD;
		16'hB4BE: out_word = 8'h20;
		16'hB4BF: out_word = 8'h1F;
		16'hB4C0: out_word = 8'hCD;
		16'hB4C1: out_word = 8'hF6;
		16'hB4C2: out_word = 8'h34;
		16'hB4C3: out_word = 8'h30;
		16'hB4C4: out_word = 8'hCC;
		16'hB4C5: out_word = 8'hEB;
		16'hB4C6: out_word = 8'h7D;
		16'hB4C7: out_word = 8'hB4;
		16'hB4C8: out_word = 8'h37;
		16'hB4C9: out_word = 8'hC2;
		16'hB4CA: out_word = 8'h4D;
		16'hB4CB: out_word = 8'h34;
		16'hB4CC: out_word = 8'h3F;
		16'hB4CD: out_word = 8'h18;
		16'hB4CE: out_word = 8'hC2;
		16'hB4CF: out_word = 8'hE5;
		16'hB4D0: out_word = 8'h23;
		16'hB4D1: out_word = 8'h23;
		16'hB4D2: out_word = 8'h5E;
		16'hB4D3: out_word = 8'h23;
		16'hB4D4: out_word = 8'h56;
		16'hB4D5: out_word = 8'h23;
		16'hB4D6: out_word = 8'h19;
		16'hB4D7: out_word = 8'hD1;
		16'hB4D8: out_word = 8'hC9;
		16'hB4D9: out_word = 8'h7E;
		16'hB4DA: out_word = 8'hE6;
		16'hB4DB: out_word = 8'hC0;
		16'hB4DC: out_word = 8'h37;
		16'hB4DD: out_word = 8'hC8;
		16'hB4DE: out_word = 8'h3F;
		16'hB4DF: out_word = 8'hC9;
		16'hB4E0: out_word = 8'h78;
		16'hB4E1: out_word = 8'hBE;
		16'hB4E2: out_word = 8'hC0;
		16'hB4E3: out_word = 8'h79;
		16'hB4E4: out_word = 8'h23;
		16'hB4E5: out_word = 8'hBE;
		16'hB4E6: out_word = 8'h2B;
		16'hB4E7: out_word = 8'hC0;
		16'hB4E8: out_word = 8'h37;
		16'hB4E9: out_word = 8'hC9;
		16'hB4EA: out_word = 8'hE5;
		16'hB4EB: out_word = 8'h21;
		16'hB4EC: out_word = 8'h00;
		16'hB4ED: out_word = 8'h00;
		16'hB4EE: out_word = 8'h22;
		16'hB4EF: out_word = 8'hA1;
		16'hB4F0: out_word = 8'hFC;
		16'hB4F1: out_word = 8'h22;
		16'hB4F2: out_word = 8'h9F;
		16'hB4F3: out_word = 8'hFC;
		16'hB4F4: out_word = 8'hE1;
		16'hB4F5: out_word = 8'hC9;
		16'hB4F6: out_word = 8'hE5;
		16'hB4F7: out_word = 8'hC1;
		16'hB4F8: out_word = 8'h11;
		16'hB4F9: out_word = 8'h00;
		16'hB4FA: out_word = 8'h00;
		16'hB4FB: out_word = 8'h2A;
		16'hB4FC: out_word = 8'h53;
		16'hB4FD: out_word = 8'h5C;
		16'hB4FE: out_word = 8'hCD;
		16'hB4FF: out_word = 8'hD9;
		16'hB500: out_word = 8'h34;
		16'hB501: out_word = 8'hD0;
		16'hB502: out_word = 8'hCD;
		16'hB503: out_word = 8'hE0;
		16'hB504: out_word = 8'h34;
		16'hB505: out_word = 8'hD8;
		16'hB506: out_word = 8'h78;
		16'hB507: out_word = 8'hB1;
		16'hB508: out_word = 8'h37;
		16'hB509: out_word = 8'hC8;
		16'hB50A: out_word = 8'hCD;
		16'hB50B: out_word = 8'hCF;
		16'hB50C: out_word = 8'h34;
		16'hB50D: out_word = 8'hCD;
		16'hB50E: out_word = 8'hD9;
		16'hB50F: out_word = 8'h34;
		16'hB510: out_word = 8'hD0;
		16'hB511: out_word = 8'hCD;
		16'hB512: out_word = 8'hE0;
		16'hB513: out_word = 8'h34;
		16'hB514: out_word = 8'h30;
		16'hB515: out_word = 8'hF4;
		16'hB516: out_word = 8'hC9;
		16'hB517: out_word = 8'h2A;
		16'hB518: out_word = 8'hA1;
		16'hB519: out_word = 8'hFC;
		16'hB51A: out_word = 8'h7D;
		16'hB51B: out_word = 8'hB4;
		16'hB51C: out_word = 8'h28;
		16'hB51D: out_word = 8'h1E;
		16'hB51E: out_word = 8'h7E;
		16'hB51F: out_word = 8'h23;
		16'hB520: out_word = 8'hFE;
		16'hB521: out_word = 8'hA0;
		16'hB522: out_word = 8'h47;
		16'hB523: out_word = 8'h3E;
		16'hB524: out_word = 8'h00;
		16'hB525: out_word = 8'h20;
		16'hB526: out_word = 8'h02;
		16'hB527: out_word = 8'h3E;
		16'hB528: out_word = 8'hFF;
		16'hB529: out_word = 8'h32;
		16'hB52A: out_word = 8'h9E;
		16'hB52B: out_word = 8'hFC;
		16'hB52C: out_word = 8'h78;
		16'hB52D: out_word = 8'hCB;
		16'hB52E: out_word = 8'h7F;
		16'hB52F: out_word = 8'h28;
		16'hB530: out_word = 8'h03;
		16'hB531: out_word = 8'h21;
		16'hB532: out_word = 8'h00;
		16'hB533: out_word = 8'h00;
		16'hB534: out_word = 8'h22;
		16'hB535: out_word = 8'hA1;
		16'hB536: out_word = 8'hFC;
		16'hB537: out_word = 8'hE6;
		16'hB538: out_word = 8'h7F;
		16'hB539: out_word = 8'hC3;
		16'hB53A: out_word = 8'h8F;
		16'hB53B: out_word = 8'h35;
		16'hB53C: out_word = 8'h2A;
		16'hB53D: out_word = 8'h9F;
		16'hB53E: out_word = 8'hFC;
		16'hB53F: out_word = 8'h7D;
		16'hB540: out_word = 8'hB4;
		16'hB541: out_word = 8'hCA;
		16'hB542: out_word = 8'h91;
		16'hB543: out_word = 8'h35;
		16'hB544: out_word = 8'hCD;
		16'hB545: out_word = 8'h20;
		16'hB546: out_word = 8'h1F;
		16'hB547: out_word = 8'h7E;
		16'hB548: out_word = 8'hFE;
		16'hB549: out_word = 8'h0E;
		16'hB54A: out_word = 8'h20;
		16'hB54B: out_word = 8'h08;
		16'hB54C: out_word = 8'h23;
		16'hB54D: out_word = 8'h23;
		16'hB54E: out_word = 8'h23;
		16'hB54F: out_word = 8'h23;
		16'hB550: out_word = 8'h23;
		16'hB551: out_word = 8'h23;
		16'hB552: out_word = 8'h18;
		16'hB553: out_word = 8'hF3;
		16'hB554: out_word = 8'hCD;
		16'hB555: out_word = 8'h45;
		16'hB556: out_word = 8'h1F;
		16'hB557: out_word = 8'h23;
		16'hB558: out_word = 8'h22;
		16'hB559: out_word = 8'h9F;
		16'hB55A: out_word = 8'hFC;
		16'hB55B: out_word = 8'hFE;
		16'hB55C: out_word = 8'hA5;
		16'hB55D: out_word = 8'h38;
		16'hB55E: out_word = 8'h08;
		16'hB55F: out_word = 8'hD6;
		16'hB560: out_word = 8'hA5;
		16'hB561: out_word = 8'hCD;
		16'hB562: out_word = 8'hAE;
		16'hB563: out_word = 8'hFC;
		16'hB564: out_word = 8'hC3;
		16'hB565: out_word = 8'h17;
		16'hB566: out_word = 8'h35;
		16'hB567: out_word = 8'hFE;
		16'hB568: out_word = 8'hA3;
		16'hB569: out_word = 8'h38;
		16'hB56A: out_word = 8'h10;
		16'hB56B: out_word = 8'h20;
		16'hB56C: out_word = 8'h05;
		16'hB56D: out_word = 8'h21;
		16'hB56E: out_word = 8'h94;
		16'hB56F: out_word = 8'h35;
		16'hB570: out_word = 8'h18;
		16'hB571: out_word = 8'h03;
		16'hB572: out_word = 8'h21;
		16'hB573: out_word = 8'h9C;
		16'hB574: out_word = 8'h35;
		16'hB575: out_word = 8'hCD;
		16'hB576: out_word = 8'hFD;
		16'hB577: out_word = 8'hFC;
		16'hB578: out_word = 8'hC3;
		16'hB579: out_word = 8'h17;
		16'hB57A: out_word = 8'h35;
		16'hB57B: out_word = 8'hF5;
		16'hB57C: out_word = 8'h3E;
		16'hB57D: out_word = 8'h00;
		16'hB57E: out_word = 8'h32;
		16'hB57F: out_word = 8'h9E;
		16'hB580: out_word = 8'hFC;
		16'hB581: out_word = 8'hF1;
		16'hB582: out_word = 8'hFE;
		16'hB583: out_word = 8'h0D;
		16'hB584: out_word = 8'h20;
		16'hB585: out_word = 8'h09;
		16'hB586: out_word = 8'h21;
		16'hB587: out_word = 8'h00;
		16'hB588: out_word = 8'h00;
		16'hB589: out_word = 8'h22;
		16'hB58A: out_word = 8'hA1;
		16'hB58B: out_word = 8'hFC;
		16'hB58C: out_word = 8'h22;
		16'hB58D: out_word = 8'h9F;
		16'hB58E: out_word = 8'hFC;
		16'hB58F: out_word = 8'h37;
		16'hB590: out_word = 8'hC9;
		16'hB591: out_word = 8'h37;
		16'hB592: out_word = 8'h3F;
		16'hB593: out_word = 8'hC9;
		16'hB594: out_word = 8'h53;
		16'hB595: out_word = 8'h50;
		16'hB596: out_word = 8'h45;
		16'hB597: out_word = 8'h43;
		16'hB598: out_word = 8'h54;
		16'hB599: out_word = 8'h52;
		16'hB59A: out_word = 8'h55;
		16'hB59B: out_word = 8'hCD;
		16'hB59C: out_word = 8'h50;
		16'hB59D: out_word = 8'h4C;
		16'hB59E: out_word = 8'h41;
		16'hB59F: out_word = 8'hD9;
		16'hB5A0: out_word = 8'h47;
		16'hB5A1: out_word = 8'h4F;
		16'hB5A2: out_word = 8'h54;
		16'hB5A3: out_word = 8'hCF;
		16'hB5A4: out_word = 8'h47;
		16'hB5A5: out_word = 8'h4F;
		16'hB5A6: out_word = 8'h53;
		16'hB5A7: out_word = 8'h55;
		16'hB5A8: out_word = 8'hC2;
		16'hB5A9: out_word = 8'h44;
		16'hB5AA: out_word = 8'h45;
		16'hB5AB: out_word = 8'h46;
		16'hB5AC: out_word = 8'h46;
		16'hB5AD: out_word = 8'hCE;
		16'hB5AE: out_word = 8'h4F;
		16'hB5AF: out_word = 8'h50;
		16'hB5B0: out_word = 8'h45;
		16'hB5B1: out_word = 8'h4E;
		16'hB5B2: out_word = 8'hA3;
		16'hB5B3: out_word = 8'h43;
		16'hB5B4: out_word = 8'h4C;
		16'hB5B5: out_word = 8'h4F;
		16'hB5B6: out_word = 8'h53;
		16'hB5B7: out_word = 8'h45;
		16'hB5B8: out_word = 8'hA3;
		16'hB5B9: out_word = 8'h02;
		16'hB5BA: out_word = 8'h01;
		16'hB5BB: out_word = 8'h05;
		16'hB5BC: out_word = 8'h21;
		16'hB5BD: out_word = 8'hB9;
		16'hB5BE: out_word = 8'h35;
		16'hB5BF: out_word = 8'h11;
		16'hB5C0: out_word = 8'h6A;
		16'hB5C1: out_word = 8'hFD;
		16'hB5C2: out_word = 8'hC3;
		16'hB5C3: out_word = 8'hBA;
		16'hB5C4: out_word = 8'h3F;
		16'hB5C5: out_word = 8'h68;
		16'hB5C6: out_word = 8'h26;
		16'hB5C7: out_word = 8'h00;
		16'hB5C8: out_word = 8'h19;
		16'hB5C9: out_word = 8'h77;
		16'hB5CA: out_word = 8'h04;
		16'hB5CB: out_word = 8'hC9;
		16'hB5CC: out_word = 8'hCD;
		16'hB5CD: out_word = 8'hE6;
		16'hB5CE: out_word = 8'h35;
		16'hB5CF: out_word = 8'h7E;
		16'hB5D0: out_word = 8'hF6;
		16'hB5D1: out_word = 8'h18;
		16'hB5D2: out_word = 8'h77;
		16'hB5D3: out_word = 8'h21;
		16'hB5D4: out_word = 8'h6A;
		16'hB5D5: out_word = 8'hFD;
		16'hB5D6: out_word = 8'hCB;
		16'hB5D7: out_word = 8'hC6;
		16'hB5D8: out_word = 8'h37;
		16'hB5D9: out_word = 8'hC9;
		16'hB5DA: out_word = 8'hCD;
		16'hB5DB: out_word = 8'hE6;
		16'hB5DC: out_word = 8'h35;
		16'hB5DD: out_word = 8'hCB;
		16'hB5DE: out_word = 8'hDE;
		16'hB5DF: out_word = 8'h21;
		16'hB5E0: out_word = 8'h6A;
		16'hB5E1: out_word = 8'hFD;
		16'hB5E2: out_word = 8'hCB;
		16'hB5E3: out_word = 8'hC6;
		16'hB5E4: out_word = 8'h37;
		16'hB5E5: out_word = 8'hC9;
		16'hB5E6: out_word = 8'h68;
		16'hB5E7: out_word = 8'h26;
		16'hB5E8: out_word = 8'h00;
		16'hB5E9: out_word = 8'h19;
		16'hB5EA: out_word = 8'h3E;
		16'hB5EB: out_word = 8'h20;
		16'hB5EC: out_word = 8'hB8;
		16'hB5ED: out_word = 8'hC8;
		16'hB5EE: out_word = 8'h36;
		16'hB5EF: out_word = 8'h00;
		16'hB5F0: out_word = 8'h23;
		16'hB5F1: out_word = 8'h04;
		16'hB5F2: out_word = 8'h18;
		16'hB5F3: out_word = 8'hF8;
		16'hB5F4: out_word = 8'h3A;
		16'hB5F5: out_word = 8'h6B;
		16'hB5F6: out_word = 8'hFD;
		16'hB5F7: out_word = 8'h06;
		16'hB5F8: out_word = 8'h00;
		16'hB5F9: out_word = 8'h26;
		16'hB5FA: out_word = 8'h00;
		16'hB5FB: out_word = 8'h68;
		16'hB5FC: out_word = 8'h19;
		16'hB5FD: out_word = 8'h36;
		16'hB5FE: out_word = 8'h00;
		16'hB5FF: out_word = 8'h04;
		16'hB600: out_word = 8'h3D;
		16'hB601: out_word = 8'h20;
		16'hB602: out_word = 8'hF6;
		16'hB603: out_word = 8'hC9;
		16'hB604: out_word = 8'hC5;
		16'hB605: out_word = 8'hD5;
		16'hB606: out_word = 8'hE5;
		16'hB607: out_word = 8'hE5;
		16'hB608: out_word = 8'h21;
		16'hB609: out_word = 8'hF5;
		16'hB60A: out_word = 8'hEE;
		16'hB60B: out_word = 8'hCB;
		16'hB60C: out_word = 8'h56;
		16'hB60D: out_word = 8'hE1;
		16'hB60E: out_word = 8'h20;
		16'hB60F: out_word = 8'h04;
		16'hB610: out_word = 8'h41;
		16'hB611: out_word = 8'hCD;
		16'hB612: out_word = 8'h1E;
		16'hB613: out_word = 8'h3B;
		16'hB614: out_word = 8'hE1;
		16'hB615: out_word = 8'hD1;
		16'hB616: out_word = 8'hC1;
		16'hB617: out_word = 8'hC9;
		16'hB618: out_word = 8'hC5;
		16'hB619: out_word = 8'hD5;
		16'hB61A: out_word = 8'hE5;
		16'hB61B: out_word = 8'hE5;
		16'hB61C: out_word = 8'h21;
		16'hB61D: out_word = 8'hF5;
		16'hB61E: out_word = 8'hEE;
		16'hB61F: out_word = 8'hCB;
		16'hB620: out_word = 8'h56;
		16'hB621: out_word = 8'hE1;
		16'hB622: out_word = 8'h20;
		16'hB623: out_word = 8'h04;
		16'hB624: out_word = 8'h59;
		16'hB625: out_word = 8'hCD;
		16'hB626: out_word = 8'hBF;
		16'hB627: out_word = 8'h3A;
		16'hB628: out_word = 8'hE1;
		16'hB629: out_word = 8'hD1;
		16'hB62A: out_word = 8'hC1;
		16'hB62B: out_word = 8'hC9;
		16'hB62C: out_word = 8'hC5;
		16'hB62D: out_word = 8'hD5;
		16'hB62E: out_word = 8'hE5;
		16'hB62F: out_word = 8'hE5;
		16'hB630: out_word = 8'h21;
		16'hB631: out_word = 8'hF5;
		16'hB632: out_word = 8'hEE;
		16'hB633: out_word = 8'hCB;
		16'hB634: out_word = 8'h56;
		16'hB635: out_word = 8'hE1;
		16'hB636: out_word = 8'h20;
		16'hB637: out_word = 8'h04;
		16'hB638: out_word = 8'h59;
		16'hB639: out_word = 8'hCD;
		16'hB63A: out_word = 8'hC6;
		16'hB63B: out_word = 8'h3A;
		16'hB63C: out_word = 8'hE1;
		16'hB63D: out_word = 8'hD1;
		16'hB63E: out_word = 8'hC1;
		16'hB63F: out_word = 8'hC9;
		16'hB640: out_word = 8'hF5;
		16'hB641: out_word = 8'hC5;
		16'hB642: out_word = 8'hD5;
		16'hB643: out_word = 8'hE5;
		16'hB644: out_word = 8'h78;
		16'hB645: out_word = 8'h41;
		16'hB646: out_word = 8'h4F;
		16'hB647: out_word = 8'hCD;
		16'hB648: out_word = 8'h9D;
		16'hB649: out_word = 8'h3A;
		16'hB64A: out_word = 8'hE1;
		16'hB64B: out_word = 8'hD1;
		16'hB64C: out_word = 8'hC1;
		16'hB64D: out_word = 8'hF1;
		16'hB64E: out_word = 8'hC9;
		16'hB64F: out_word = 8'hF5;
		16'hB650: out_word = 8'hC5;
		16'hB651: out_word = 8'hD5;
		16'hB652: out_word = 8'hE5;
		16'hB653: out_word = 8'h78;
		16'hB654: out_word = 8'h41;
		16'hB655: out_word = 8'h4F;
		16'hB656: out_word = 8'hCD;
		16'hB657: out_word = 8'hB2;
		16'hB658: out_word = 8'h3A;
		16'hB659: out_word = 8'hE1;
		16'hB65A: out_word = 8'hD1;
		16'hB65B: out_word = 8'hC1;
		16'hB65C: out_word = 8'hF1;
		16'hB65D: out_word = 8'hC9;
		16'hB65E: out_word = 8'h3E;
		16'hB65F: out_word = 8'h00;
		16'hB660: out_word = 8'h32;
		16'hB661: out_word = 8'h41;
		16'hB662: out_word = 8'h5C;
		16'hB663: out_word = 8'h3E;
		16'hB664: out_word = 8'h02;
		16'hB665: out_word = 8'h32;
		16'hB666: out_word = 8'h0A;
		16'hB667: out_word = 8'h5C;
		16'hB668: out_word = 8'h21;
		16'hB669: out_word = 8'h3B;
		16'hB66A: out_word = 8'h5C;
		16'hB66B: out_word = 8'h7E;
		16'hB66C: out_word = 8'hF6;
		16'hB66D: out_word = 8'h0C;
		16'hB66E: out_word = 8'h77;
		16'hB66F: out_word = 8'h21;
		16'hB670: out_word = 8'h0D;
		16'hB671: out_word = 8'hEC;
		16'hB672: out_word = 8'hCB;
		16'hB673: out_word = 8'h66;
		16'hB674: out_word = 8'h21;
		16'hB675: out_word = 8'h66;
		16'hB676: out_word = 8'h5B;
		16'hB677: out_word = 8'h20;
		16'hB678: out_word = 8'h03;
		16'hB679: out_word = 8'hCB;
		16'hB67A: out_word = 8'h86;
		16'hB67B: out_word = 8'hC9;
		16'hB67C: out_word = 8'hCB;
		16'hB67D: out_word = 8'hC6;
		16'hB67E: out_word = 8'hC9;
		16'hB67F: out_word = 8'hE5;
		16'hB680: out_word = 8'h21;
		16'hB681: out_word = 8'h3B;
		16'hB682: out_word = 8'h5C;
		16'hB683: out_word = 8'hCB;
		16'hB684: out_word = 8'h6E;
		16'hB685: out_word = 8'h28;
		16'hB686: out_word = 8'hFC;
		16'hB687: out_word = 8'hCB;
		16'hB688: out_word = 8'hAE;
		16'hB689: out_word = 8'h3A;
		16'hB68A: out_word = 8'h08;
		16'hB68B: out_word = 8'h5C;
		16'hB68C: out_word = 8'h21;
		16'hB68D: out_word = 8'h41;
		16'hB68E: out_word = 8'h5C;
		16'hB68F: out_word = 8'hCB;
		16'hB690: out_word = 8'h86;
		16'hB691: out_word = 8'hFE;
		16'hB692: out_word = 8'h20;
		16'hB693: out_word = 8'h30;
		16'hB694: out_word = 8'h0D;
		16'hB695: out_word = 8'hFE;
		16'hB696: out_word = 8'h10;
		16'hB697: out_word = 8'h30;
		16'hB698: out_word = 8'hE7;
		16'hB699: out_word = 8'hFE;
		16'hB69A: out_word = 8'h06;
		16'hB69B: out_word = 8'h38;
		16'hB69C: out_word = 8'hE3;
		16'hB69D: out_word = 8'hCD;
		16'hB69E: out_word = 8'hA4;
		16'hB69F: out_word = 8'h36;
		16'hB6A0: out_word = 8'h30;
		16'hB6A1: out_word = 8'hDE;
		16'hB6A2: out_word = 8'hE1;
		16'hB6A3: out_word = 8'hC9;
		16'hB6A4: out_word = 8'hEF;
		16'hB6A5: out_word = 8'hDB;
		16'hB6A6: out_word = 8'h10;
		16'hB6A7: out_word = 8'hC9;
		16'hB6A8: out_word = 8'hE5;
		16'hB6A9: out_word = 8'hCD;
		16'hB6AA: out_word = 8'h3B;
		16'hB6AB: out_word = 8'h37;
		16'hB6AC: out_word = 8'h21;
		16'hB6AD: out_word = 8'h3C;
		16'hB6AE: out_word = 8'h5C;
		16'hB6AF: out_word = 8'hCB;
		16'hB6B0: out_word = 8'h86;
		16'hB6B1: out_word = 8'hE1;
		16'hB6B2: out_word = 8'h5E;
		16'hB6B3: out_word = 8'h23;
		16'hB6B4: out_word = 8'hE5;
		16'hB6B5: out_word = 8'h21;
		16'hB6B6: out_word = 8'hEC;
		16'hB6B7: out_word = 8'h37;
		16'hB6B8: out_word = 8'hCD;
		16'hB6B9: out_word = 8'h33;
		16'hB6BA: out_word = 8'h37;
		16'hB6BB: out_word = 8'hE1;
		16'hB6BC: out_word = 8'hCD;
		16'hB6BD: out_word = 8'h33;
		16'hB6BE: out_word = 8'h37;
		16'hB6BF: out_word = 8'hE5;
		16'hB6C0: out_word = 8'hCD;
		16'hB6C1: out_word = 8'h22;
		16'hB6C2: out_word = 8'h38;
		16'hB6C3: out_word = 8'h21;
		16'hB6C4: out_word = 8'hFA;
		16'hB6C5: out_word = 8'h37;
		16'hB6C6: out_word = 8'hCD;
		16'hB6C7: out_word = 8'h33;
		16'hB6C8: out_word = 8'h37;
		16'hB6C9: out_word = 8'hE1;
		16'hB6CA: out_word = 8'hD5;
		16'hB6CB: out_word = 8'h01;
		16'hB6CC: out_word = 8'h07;
		16'hB6CD: out_word = 8'h08;
		16'hB6CE: out_word = 8'hCD;
		16'hB6CF: out_word = 8'h2B;
		16'hB6D0: out_word = 8'h37;
		16'hB6D1: out_word = 8'hC5;
		16'hB6D2: out_word = 8'h06;
		16'hB6D3: out_word = 8'h0C;
		16'hB6D4: out_word = 8'h3E;
		16'hB6D5: out_word = 8'h20;
		16'hB6D6: out_word = 8'hD7;
		16'hB6D7: out_word = 8'h7E;
		16'hB6D8: out_word = 8'h23;
		16'hB6D9: out_word = 8'hFE;
		16'hB6DA: out_word = 8'h80;
		16'hB6DB: out_word = 8'h30;
		16'hB6DC: out_word = 8'h03;
		16'hB6DD: out_word = 8'hD7;
		16'hB6DE: out_word = 8'h10;
		16'hB6DF: out_word = 8'hF7;
		16'hB6E0: out_word = 8'hE6;
		16'hB6E1: out_word = 8'h7F;
		16'hB6E2: out_word = 8'hD7;
		16'hB6E3: out_word = 8'h3E;
		16'hB6E4: out_word = 8'h20;
		16'hB6E5: out_word = 8'hD7;
		16'hB6E6: out_word = 8'h10;
		16'hB6E7: out_word = 8'hFB;
		16'hB6E8: out_word = 8'hC1;
		16'hB6E9: out_word = 8'h04;
		16'hB6EA: out_word = 8'hCD;
		16'hB6EB: out_word = 8'h2B;
		16'hB6EC: out_word = 8'h37;
		16'hB6ED: out_word = 8'h1D;
		16'hB6EE: out_word = 8'h20;
		16'hB6EF: out_word = 8'hE1;
		16'hB6F0: out_word = 8'h21;
		16'hB6F1: out_word = 8'h38;
		16'hB6F2: out_word = 8'h6F;
		16'hB6F3: out_word = 8'hD1;
		16'hB6F4: out_word = 8'hCB;
		16'hB6F5: out_word = 8'h23;
		16'hB6F6: out_word = 8'hCB;
		16'hB6F7: out_word = 8'h23;
		16'hB6F8: out_word = 8'hCB;
		16'hB6F9: out_word = 8'h23;
		16'hB6FA: out_word = 8'h53;
		16'hB6FB: out_word = 8'h15;
		16'hB6FC: out_word = 8'h1E;
		16'hB6FD: out_word = 8'h6F;
		16'hB6FE: out_word = 8'h01;
		16'hB6FF: out_word = 8'h00;
		16'hB700: out_word = 8'hFF;
		16'hB701: out_word = 8'h7A;
		16'hB702: out_word = 8'hCD;
		16'hB703: out_word = 8'h19;
		16'hB704: out_word = 8'h37;
		16'hB705: out_word = 8'h01;
		16'hB706: out_word = 8'h01;
		16'hB707: out_word = 8'h00;
		16'hB708: out_word = 8'h7B;
		16'hB709: out_word = 8'hCD;
		16'hB70A: out_word = 8'h19;
		16'hB70B: out_word = 8'h37;
		16'hB70C: out_word = 8'h01;
		16'hB70D: out_word = 8'h00;
		16'hB70E: out_word = 8'h01;
		16'hB70F: out_word = 8'h7A;
		16'hB710: out_word = 8'h3C;
		16'hB711: out_word = 8'hCD;
		16'hB712: out_word = 8'h19;
		16'hB713: out_word = 8'h37;
		16'hB714: out_word = 8'hAF;
		16'hB715: out_word = 8'hCD;
		16'hB716: out_word = 8'hCA;
		16'hB717: out_word = 8'h37;
		16'hB718: out_word = 8'hC9;
		16'hB719: out_word = 8'hF5;
		16'hB71A: out_word = 8'hE5;
		16'hB71B: out_word = 8'hD5;
		16'hB71C: out_word = 8'hC5;
		16'hB71D: out_word = 8'h44;
		16'hB71E: out_word = 8'h4D;
		16'hB71F: out_word = 8'hEF;
		16'hB720: out_word = 8'hE9;
		16'hB721: out_word = 8'h22;
		16'hB722: out_word = 8'hC1;
		16'hB723: out_word = 8'hD1;
		16'hB724: out_word = 8'hE1;
		16'hB725: out_word = 8'hF1;
		16'hB726: out_word = 8'h09;
		16'hB727: out_word = 8'h3D;
		16'hB728: out_word = 8'h20;
		16'hB729: out_word = 8'hEF;
		16'hB72A: out_word = 8'hC9;
		16'hB72B: out_word = 8'h3E;
		16'hB72C: out_word = 8'h16;
		16'hB72D: out_word = 8'hD7;
		16'hB72E: out_word = 8'h78;
		16'hB72F: out_word = 8'hD7;
		16'hB730: out_word = 8'h79;
		16'hB731: out_word = 8'hD7;
		16'hB732: out_word = 8'hC9;
		16'hB733: out_word = 8'h7E;
		16'hB734: out_word = 8'h23;
		16'hB735: out_word = 8'hFE;
		16'hB736: out_word = 8'hFF;
		16'hB737: out_word = 8'hC8;
		16'hB738: out_word = 8'hD7;
		16'hB739: out_word = 8'h18;
		16'hB73A: out_word = 8'hF8;
		16'hB73B: out_word = 8'h37;
		16'hB73C: out_word = 8'h18;
		16'hB73D: out_word = 8'h01;
		16'hB73E: out_word = 8'hA7;
		16'hB73F: out_word = 8'h11;
		16'hB740: out_word = 8'hF6;
		16'hB741: out_word = 8'hEE;
		16'hB742: out_word = 8'h21;
		16'hB743: out_word = 8'h3C;
		16'hB744: out_word = 8'h5C;
		16'hB745: out_word = 8'h38;
		16'hB746: out_word = 8'h01;
		16'hB747: out_word = 8'hEB;
		16'hB748: out_word = 8'hED;
		16'hB749: out_word = 8'hA0;
		16'hB74A: out_word = 8'h38;
		16'hB74B: out_word = 8'h01;
		16'hB74C: out_word = 8'hEB;
		16'hB74D: out_word = 8'h21;
		16'hB74E: out_word = 8'h7D;
		16'hB74F: out_word = 8'h5C;
		16'hB750: out_word = 8'h38;
		16'hB751: out_word = 8'h01;
		16'hB752: out_word = 8'hEB;
		16'hB753: out_word = 8'h01;
		16'hB754: out_word = 8'h14;
		16'hB755: out_word = 8'h00;
		16'hB756: out_word = 8'hED;
		16'hB757: out_word = 8'hB0;
		16'hB758: out_word = 8'h38;
		16'hB759: out_word = 8'h01;
		16'hB75A: out_word = 8'hEB;
		16'hB75B: out_word = 8'h08;
		16'hB75C: out_word = 8'h01;
		16'hB75D: out_word = 8'h07;
		16'hB75E: out_word = 8'h07;
		16'hB75F: out_word = 8'hCD;
		16'hB760: out_word = 8'h94;
		16'hB761: out_word = 8'h3B;
		16'hB762: out_word = 8'hDD;
		16'hB763: out_word = 8'h7E;
		16'hB764: out_word = 8'h01;
		16'hB765: out_word = 8'h80;
		16'hB766: out_word = 8'h47;
		16'hB767: out_word = 8'h3E;
		16'hB768: out_word = 8'h0C;
		16'hB769: out_word = 8'hC5;
		16'hB76A: out_word = 8'hF5;
		16'hB76B: out_word = 8'hD5;
		16'hB76C: out_word = 8'hEF;
		16'hB76D: out_word = 8'h9B;
		16'hB76E: out_word = 8'h0E;
		16'hB76F: out_word = 8'h01;
		16'hB770: out_word = 8'h07;
		16'hB771: out_word = 8'h00;
		16'hB772: out_word = 8'h09;
		16'hB773: out_word = 8'hD1;
		16'hB774: out_word = 8'hCD;
		16'hB775: out_word = 8'h7E;
		16'hB776: out_word = 8'h37;
		16'hB777: out_word = 8'hF1;
		16'hB778: out_word = 8'hC1;
		16'hB779: out_word = 8'h05;
		16'hB77A: out_word = 8'h3D;
		16'hB77B: out_word = 8'h20;
		16'hB77C: out_word = 8'hEC;
		16'hB77D: out_word = 8'hC9;
		16'hB77E: out_word = 8'h01;
		16'hB77F: out_word = 8'h0E;
		16'hB780: out_word = 8'h08;
		16'hB781: out_word = 8'hC5;
		16'hB782: out_word = 8'h06;
		16'hB783: out_word = 8'h00;
		16'hB784: out_word = 8'hE5;
		16'hB785: out_word = 8'h08;
		16'hB786: out_word = 8'h38;
		16'hB787: out_word = 8'h01;
		16'hB788: out_word = 8'hEB;
		16'hB789: out_word = 8'hED;
		16'hB78A: out_word = 8'hB0;
		16'hB78B: out_word = 8'h38;
		16'hB78C: out_word = 8'h01;
		16'hB78D: out_word = 8'hEB;
		16'hB78E: out_word = 8'h08;
		16'hB78F: out_word = 8'hE1;
		16'hB790: out_word = 8'h24;
		16'hB791: out_word = 8'hC1;
		16'hB792: out_word = 8'h10;
		16'hB793: out_word = 8'hED;
		16'hB794: out_word = 8'hC5;
		16'hB795: out_word = 8'hD5;
		16'hB796: out_word = 8'hEF;
		16'hB797: out_word = 8'h88;
		16'hB798: out_word = 8'h0E;
		16'hB799: out_word = 8'hEB;
		16'hB79A: out_word = 8'hD1;
		16'hB79B: out_word = 8'hC1;
		16'hB79C: out_word = 8'h08;
		16'hB79D: out_word = 8'h38;
		16'hB79E: out_word = 8'h01;
		16'hB79F: out_word = 8'hEB;
		16'hB7A0: out_word = 8'hED;
		16'hB7A1: out_word = 8'hB0;
		16'hB7A2: out_word = 8'h38;
		16'hB7A3: out_word = 8'h01;
		16'hB7A4: out_word = 8'hEB;
		16'hB7A5: out_word = 8'h08;
		16'hB7A6: out_word = 8'hC9;
		16'hB7A7: out_word = 8'hCD;
		16'hB7A8: out_word = 8'hCA;
		16'hB7A9: out_word = 8'h37;
		16'hB7AA: out_word = 8'h3D;
		16'hB7AB: out_word = 8'hF2;
		16'hB7AC: out_word = 8'hB1;
		16'hB7AD: out_word = 8'h37;
		16'hB7AE: out_word = 8'h7E;
		16'hB7AF: out_word = 8'h3D;
		16'hB7B0: out_word = 8'h3D;
		16'hB7B1: out_word = 8'hCD;
		16'hB7B2: out_word = 8'hCA;
		16'hB7B3: out_word = 8'h37;
		16'hB7B4: out_word = 8'h37;
		16'hB7B5: out_word = 8'hC9;
		16'hB7B6: out_word = 8'hD5;
		16'hB7B7: out_word = 8'hCD;
		16'hB7B8: out_word = 8'hCA;
		16'hB7B9: out_word = 8'h37;
		16'hB7BA: out_word = 8'h3C;
		16'hB7BB: out_word = 8'h57;
		16'hB7BC: out_word = 8'h7E;
		16'hB7BD: out_word = 8'h3D;
		16'hB7BE: out_word = 8'h3D;
		16'hB7BF: out_word = 8'hBA;
		16'hB7C0: out_word = 8'h7A;
		16'hB7C1: out_word = 8'hF2;
		16'hB7C2: out_word = 8'hC5;
		16'hB7C3: out_word = 8'h37;
		16'hB7C4: out_word = 8'hAF;
		16'hB7C5: out_word = 8'hCD;
		16'hB7C6: out_word = 8'hCA;
		16'hB7C7: out_word = 8'h37;
		16'hB7C8: out_word = 8'hD1;
		16'hB7C9: out_word = 8'hC9;
		16'hB7CA: out_word = 8'hF5;
		16'hB7CB: out_word = 8'hE5;
		16'hB7CC: out_word = 8'hD5;
		16'hB7CD: out_word = 8'h21;
		16'hB7CE: out_word = 8'h07;
		16'hB7CF: out_word = 8'h59;
		16'hB7D0: out_word = 8'h11;
		16'hB7D1: out_word = 8'h20;
		16'hB7D2: out_word = 8'h00;
		16'hB7D3: out_word = 8'hA7;
		16'hB7D4: out_word = 8'h28;
		16'hB7D5: out_word = 8'h04;
		16'hB7D6: out_word = 8'h19;
		16'hB7D7: out_word = 8'h3D;
		16'hB7D8: out_word = 8'h20;
		16'hB7D9: out_word = 8'hFC;
		16'hB7DA: out_word = 8'h3E;
		16'hB7DB: out_word = 8'h78;
		16'hB7DC: out_word = 8'hBE;
		16'hB7DD: out_word = 8'h20;
		16'hB7DE: out_word = 8'h02;
		16'hB7DF: out_word = 8'h3E;
		16'hB7E0: out_word = 8'h68;
		16'hB7E1: out_word = 8'h16;
		16'hB7E2: out_word = 8'h0E;
		16'hB7E3: out_word = 8'h77;
		16'hB7E4: out_word = 8'h23;
		16'hB7E5: out_word = 8'h15;
		16'hB7E6: out_word = 8'h20;
		16'hB7E7: out_word = 8'hFB;
		16'hB7E8: out_word = 8'hD1;
		16'hB7E9: out_word = 8'hE1;
		16'hB7EA: out_word = 8'hF1;
		16'hB7EB: out_word = 8'hC9;
		16'hB7EC: out_word = 8'h16;
		16'hB7ED: out_word = 8'h07;
		16'hB7EE: out_word = 8'h07;
		16'hB7EF: out_word = 8'h15;
		16'hB7F0: out_word = 8'h00;
		16'hB7F1: out_word = 8'h14;
		16'hB7F2: out_word = 8'h00;
		16'hB7F3: out_word = 8'h10;
		16'hB7F4: out_word = 8'h07;
		16'hB7F5: out_word = 8'h11;
		16'hB7F6: out_word = 8'h00;
		16'hB7F7: out_word = 8'h13;
		16'hB7F8: out_word = 8'h01;
		16'hB7F9: out_word = 8'hFF;
		16'hB7FA: out_word = 8'h11;
		16'hB7FB: out_word = 8'h00;
		16'hB7FC: out_word = 8'h20;
		16'hB7FD: out_word = 8'h11;
		16'hB7FE: out_word = 8'h07;
		16'hB7FF: out_word = 8'h10;
		16'hB800: out_word = 8'h00;
		16'hB801: out_word = 8'hFF;
		16'hB802: out_word = 8'h01;
		16'hB803: out_word = 8'h03;
		16'hB804: out_word = 8'h07;
		16'hB805: out_word = 8'h0F;
		16'hB806: out_word = 8'h1F;
		16'hB807: out_word = 8'h3F;
		16'hB808: out_word = 8'h7F;
		16'hB809: out_word = 8'hFF;
		16'hB80A: out_word = 8'hFE;
		16'hB80B: out_word = 8'hFC;
		16'hB80C: out_word = 8'hF8;
		16'hB80D: out_word = 8'hF0;
		16'hB80E: out_word = 8'hE0;
		16'hB80F: out_word = 8'hC0;
		16'hB810: out_word = 8'h80;
		16'hB811: out_word = 8'h00;
		16'hB812: out_word = 8'h10;
		16'hB813: out_word = 8'h02;
		16'hB814: out_word = 8'h20;
		16'hB815: out_word = 8'h11;
		16'hB816: out_word = 8'h06;
		16'hB817: out_word = 8'h21;
		16'hB818: out_word = 8'h10;
		16'hB819: out_word = 8'h04;
		16'hB81A: out_word = 8'h20;
		16'hB81B: out_word = 8'h11;
		16'hB81C: out_word = 8'h05;
		16'hB81D: out_word = 8'h21;
		16'hB81E: out_word = 8'h10;
		16'hB81F: out_word = 8'h00;
		16'hB820: out_word = 8'h20;
		16'hB821: out_word = 8'hFF;
		16'hB822: out_word = 8'hC5;
		16'hB823: out_word = 8'hD5;
		16'hB824: out_word = 8'hE5;
		16'hB825: out_word = 8'h21;
		16'hB826: out_word = 8'h02;
		16'hB827: out_word = 8'h38;
		16'hB828: out_word = 8'h11;
		16'hB829: out_word = 8'h98;
		16'hB82A: out_word = 8'h5B;
		16'hB82B: out_word = 8'h01;
		16'hB82C: out_word = 8'h10;
		16'hB82D: out_word = 8'h00;
		16'hB82E: out_word = 8'hED;
		16'hB82F: out_word = 8'hB0;
		16'hB830: out_word = 8'h2A;
		16'hB831: out_word = 8'h36;
		16'hB832: out_word = 8'h5C;
		16'hB833: out_word = 8'hE5;
		16'hB834: out_word = 8'h21;
		16'hB835: out_word = 8'h98;
		16'hB836: out_word = 8'h5A;
		16'hB837: out_word = 8'h22;
		16'hB838: out_word = 8'h36;
		16'hB839: out_word = 8'h5C;
		16'hB83A: out_word = 8'h21;
		16'hB83B: out_word = 8'h12;
		16'hB83C: out_word = 8'h38;
		16'hB83D: out_word = 8'hCD;
		16'hB83E: out_word = 8'h33;
		16'hB83F: out_word = 8'h37;
		16'hB840: out_word = 8'hE1;
		16'hB841: out_word = 8'h22;
		16'hB842: out_word = 8'h36;
		16'hB843: out_word = 8'h5C;
		16'hB844: out_word = 8'hE1;
		16'hB845: out_word = 8'hD1;
		16'hB846: out_word = 8'hC1;
		16'hB847: out_word = 8'hC9;
		16'hB848: out_word = 8'h21;
		16'hB849: out_word = 8'h69;
		16'hB84A: out_word = 8'h27;
		16'hB84B: out_word = 8'h18;
		16'hB84C: out_word = 8'h0D;
		16'hB84D: out_word = 8'h21;
		16'hB84E: out_word = 8'h72;
		16'hB84F: out_word = 8'h27;
		16'hB850: out_word = 8'h18;
		16'hB851: out_word = 8'h08;
		16'hB852: out_word = 8'h21;
		16'hB853: out_word = 8'h5E;
		16'hB854: out_word = 8'h27;
		16'hB855: out_word = 8'h18;
		16'hB856: out_word = 8'h03;
		16'hB857: out_word = 8'h21;
		16'hB858: out_word = 8'h84;
		16'hB859: out_word = 8'h27;
		16'hB85A: out_word = 8'hE5;
		16'hB85B: out_word = 8'hCD;
		16'hB85C: out_word = 8'h81;
		16'hB85D: out_word = 8'h38;
		16'hB85E: out_word = 8'h21;
		16'hB85F: out_word = 8'hA0;
		16'hB860: out_word = 8'h5A;
		16'hB861: out_word = 8'h06;
		16'hB862: out_word = 8'h20;
		16'hB863: out_word = 8'h3E;
		16'hB864: out_word = 8'h40;
		16'hB865: out_word = 8'h77;
		16'hB866: out_word = 8'h23;
		16'hB867: out_word = 8'h10;
		16'hB868: out_word = 8'hFC;
		16'hB869: out_word = 8'h21;
		16'hB86A: out_word = 8'hEC;
		16'hB86B: out_word = 8'h37;
		16'hB86C: out_word = 8'hCD;
		16'hB86D: out_word = 8'h33;
		16'hB86E: out_word = 8'h37;
		16'hB86F: out_word = 8'h01;
		16'hB870: out_word = 8'h00;
		16'hB871: out_word = 8'h15;
		16'hB872: out_word = 8'hCD;
		16'hB873: out_word = 8'h2B;
		16'hB874: out_word = 8'h37;
		16'hB875: out_word = 8'hD1;
		16'hB876: out_word = 8'hCD;
		16'hB877: out_word = 8'h7D;
		16'hB878: out_word = 8'h05;
		16'hB879: out_word = 8'h0E;
		16'hB87A: out_word = 8'h1A;
		16'hB87B: out_word = 8'hCD;
		16'hB87C: out_word = 8'h2B;
		16'hB87D: out_word = 8'h37;
		16'hB87E: out_word = 8'hC3;
		16'hB87F: out_word = 8'h22;
		16'hB880: out_word = 8'h38;
		16'hB881: out_word = 8'h06;
		16'hB882: out_word = 8'h15;
		16'hB883: out_word = 8'h16;
		16'hB884: out_word = 8'h17;
		16'hB885: out_word = 8'hC3;
		16'hB886: out_word = 8'h5E;
		16'hB887: out_word = 8'h3B;
		16'hB888: out_word = 8'hCD;
		16'hB889: out_word = 8'h20;
		16'hB88A: out_word = 8'h1F;
		16'hB88B: out_word = 8'hCD;
		16'hB88C: out_word = 8'h05;
		16'hB88D: out_word = 8'h3A;
		16'hB88E: out_word = 8'h7A;
		16'hB88F: out_word = 8'hB3;
		16'hB890: out_word = 8'hCA;
		16'hB891: out_word = 8'hC0;
		16'hB892: out_word = 8'h39;
		16'hB893: out_word = 8'h2A;
		16'hB894: out_word = 8'h96;
		16'hB895: out_word = 8'h5B;
		16'hB896: out_word = 8'hEF;
		16'hB897: out_word = 8'hA9;
		16'hB898: out_word = 8'h30;
		16'hB899: out_word = 8'hEB;
		16'hB89A: out_word = 8'h2A;
		16'hB89B: out_word = 8'h94;
		16'hB89C: out_word = 8'h5B;
		16'hB89D: out_word = 8'h19;
		16'hB89E: out_word = 8'h11;
		16'hB89F: out_word = 8'h10;
		16'hB8A0: out_word = 8'h27;
		16'hB8A1: out_word = 8'hB7;
		16'hB8A2: out_word = 8'hED;
		16'hB8A3: out_word = 8'h52;
		16'hB8A4: out_word = 8'hD2;
		16'hB8A5: out_word = 8'hC0;
		16'hB8A6: out_word = 8'h39;
		16'hB8A7: out_word = 8'h2A;
		16'hB8A8: out_word = 8'h53;
		16'hB8A9: out_word = 8'h5C;
		16'hB8AA: out_word = 8'hEF;
		16'hB8AB: out_word = 8'hB8;
		16'hB8AC: out_word = 8'h19;
		16'hB8AD: out_word = 8'h23;
		16'hB8AE: out_word = 8'h23;
		16'hB8AF: out_word = 8'h22;
		16'hB8B0: out_word = 8'h92;
		16'hB8B1: out_word = 8'h5B;
		16'hB8B2: out_word = 8'h23;
		16'hB8B3: out_word = 8'h23;
		16'hB8B4: out_word = 8'hED;
		16'hB8B5: out_word = 8'h53;
		16'hB8B6: out_word = 8'h6B;
		16'hB8B7: out_word = 8'h5B;
		16'hB8B8: out_word = 8'h7E;
		16'hB8B9: out_word = 8'hEF;
		16'hB8BA: out_word = 8'hB6;
		16'hB8BB: out_word = 8'h18;
		16'hB8BC: out_word = 8'hFE;
		16'hB8BD: out_word = 8'h0D;
		16'hB8BE: out_word = 8'h28;
		16'hB8BF: out_word = 8'h05;
		16'hB8C0: out_word = 8'hCD;
		16'hB8C1: out_word = 8'h0E;
		16'hB8C2: out_word = 8'h39;
		16'hB8C3: out_word = 8'h18;
		16'hB8C4: out_word = 8'hF3;
		16'hB8C5: out_word = 8'hED;
		16'hB8C6: out_word = 8'h5B;
		16'hB8C7: out_word = 8'h6B;
		16'hB8C8: out_word = 8'h5B;
		16'hB8C9: out_word = 8'h2A;
		16'hB8CA: out_word = 8'h4B;
		16'hB8CB: out_word = 8'h5C;
		16'hB8CC: out_word = 8'hA7;
		16'hB8CD: out_word = 8'hED;
		16'hB8CE: out_word = 8'h52;
		16'hB8CF: out_word = 8'hEB;
		16'hB8D0: out_word = 8'h20;
		16'hB8D1: out_word = 8'hD8;
		16'hB8D2: out_word = 8'hCD;
		16'hB8D3: out_word = 8'h05;
		16'hB8D4: out_word = 8'h3A;
		16'hB8D5: out_word = 8'h42;
		16'hB8D6: out_word = 8'h4B;
		16'hB8D7: out_word = 8'h11;
		16'hB8D8: out_word = 8'h00;
		16'hB8D9: out_word = 8'h00;
		16'hB8DA: out_word = 8'h2A;
		16'hB8DB: out_word = 8'h53;
		16'hB8DC: out_word = 8'h5C;
		16'hB8DD: out_word = 8'hC5;
		16'hB8DE: out_word = 8'hD5;
		16'hB8DF: out_word = 8'hE5;
		16'hB8E0: out_word = 8'h2A;
		16'hB8E1: out_word = 8'h96;
		16'hB8E2: out_word = 8'h5B;
		16'hB8E3: out_word = 8'hEF;
		16'hB8E4: out_word = 8'hA9;
		16'hB8E5: out_word = 8'h30;
		16'hB8E6: out_word = 8'hED;
		16'hB8E7: out_word = 8'h5B;
		16'hB8E8: out_word = 8'h94;
		16'hB8E9: out_word = 8'h5B;
		16'hB8EA: out_word = 8'h19;
		16'hB8EB: out_word = 8'hEB;
		16'hB8EC: out_word = 8'hE1;
		16'hB8ED: out_word = 8'h72;
		16'hB8EE: out_word = 8'h23;
		16'hB8EF: out_word = 8'h73;
		16'hB8F0: out_word = 8'h23;
		16'hB8F1: out_word = 8'h4E;
		16'hB8F2: out_word = 8'h23;
		16'hB8F3: out_word = 8'h46;
		16'hB8F4: out_word = 8'h23;
		16'hB8F5: out_word = 8'h09;
		16'hB8F6: out_word = 8'hD1;
		16'hB8F7: out_word = 8'h13;
		16'hB8F8: out_word = 8'hC1;
		16'hB8F9: out_word = 8'h0B;
		16'hB8FA: out_word = 8'h78;
		16'hB8FB: out_word = 8'hB1;
		16'hB8FC: out_word = 8'h20;
		16'hB8FD: out_word = 8'hDF;
		16'hB8FE: out_word = 8'hCD;
		16'hB8FF: out_word = 8'h45;
		16'hB900: out_word = 8'h1F;
		16'hB901: out_word = 8'hED;
		16'hB902: out_word = 8'h43;
		16'hB903: out_word = 8'h92;
		16'hB904: out_word = 8'h5B;
		16'hB905: out_word = 8'h37;
		16'hB906: out_word = 8'hC9;
		16'hB907: out_word = 8'hCA;
		16'hB908: out_word = 8'hF0;
		16'hB909: out_word = 8'hE1;
		16'hB90A: out_word = 8'hEC;
		16'hB90B: out_word = 8'hED;
		16'hB90C: out_word = 8'hE5;
		16'hB90D: out_word = 8'hF7;
		16'hB90E: out_word = 8'h23;
		16'hB90F: out_word = 8'h22;
		16'hB910: out_word = 8'h79;
		16'hB911: out_word = 8'h5B;
		16'hB912: out_word = 8'hEB;
		16'hB913: out_word = 8'h01;
		16'hB914: out_word = 8'h07;
		16'hB915: out_word = 8'h00;
		16'hB916: out_word = 8'h21;
		16'hB917: out_word = 8'h07;
		16'hB918: out_word = 8'h39;
		16'hB919: out_word = 8'hED;
		16'hB91A: out_word = 8'hB1;
		16'hB91B: out_word = 8'hEB;
		16'hB91C: out_word = 8'hC0;
		16'hB91D: out_word = 8'h0E;
		16'hB91E: out_word = 8'h00;
		16'hB91F: out_word = 8'h7E;
		16'hB920: out_word = 8'hFE;
		16'hB921: out_word = 8'h20;
		16'hB922: out_word = 8'h28;
		16'hB923: out_word = 8'h1B;
		16'hB924: out_word = 8'hEF;
		16'hB925: out_word = 8'h1B;
		16'hB926: out_word = 8'h2D;
		16'hB927: out_word = 8'h30;
		16'hB928: out_word = 8'h16;
		16'hB929: out_word = 8'hFE;
		16'hB92A: out_word = 8'h2E;
		16'hB92B: out_word = 8'h28;
		16'hB92C: out_word = 8'h12;
		16'hB92D: out_word = 8'hFE;
		16'hB92E: out_word = 8'h0E;
		16'hB92F: out_word = 8'h28;
		16'hB930: out_word = 8'h12;
		16'hB931: out_word = 8'hF6;
		16'hB932: out_word = 8'h20;
		16'hB933: out_word = 8'hFE;
		16'hB934: out_word = 8'h65;
		16'hB935: out_word = 8'h20;
		16'hB936: out_word = 8'h04;
		16'hB937: out_word = 8'h78;
		16'hB938: out_word = 8'hB1;
		16'hB939: out_word = 8'h20;
		16'hB93A: out_word = 8'h04;
		16'hB93B: out_word = 8'h2A;
		16'hB93C: out_word = 8'h79;
		16'hB93D: out_word = 8'h5B;
		16'hB93E: out_word = 8'hC9;
		16'hB93F: out_word = 8'h03;
		16'hB940: out_word = 8'h23;
		16'hB941: out_word = 8'h18;
		16'hB942: out_word = 8'hDC;
		16'hB943: out_word = 8'hED;
		16'hB944: out_word = 8'h43;
		16'hB945: out_word = 8'h71;
		16'hB946: out_word = 8'h5B;
		16'hB947: out_word = 8'hE5;
		16'hB948: out_word = 8'hEF;
		16'hB949: out_word = 8'hB6;
		16'hB94A: out_word = 8'h18;
		16'hB94B: out_word = 8'hCD;
		16'hB94C: out_word = 8'h36;
		16'hB94D: out_word = 8'h3A;
		16'hB94E: out_word = 8'h7E;
		16'hB94F: out_word = 8'hE1;
		16'hB950: out_word = 8'hFE;
		16'hB951: out_word = 8'h3A;
		16'hB952: out_word = 8'h28;
		16'hB953: out_word = 8'h03;
		16'hB954: out_word = 8'hFE;
		16'hB955: out_word = 8'h0D;
		16'hB956: out_word = 8'hC0;
		16'hB957: out_word = 8'h23;
		16'hB958: out_word = 8'hEF;
		16'hB959: out_word = 8'hB4;
		16'hB95A: out_word = 8'h33;
		16'hB95B: out_word = 8'hEF;
		16'hB95C: out_word = 8'hA2;
		16'hB95D: out_word = 8'h2D;
		16'hB95E: out_word = 8'h60;
		16'hB95F: out_word = 8'h69;
		16'hB960: out_word = 8'hEF;
		16'hB961: out_word = 8'h6E;
		16'hB962: out_word = 8'h19;
		16'hB963: out_word = 8'h28;
		16'hB964: out_word = 8'h0A;
		16'hB965: out_word = 8'h7E;
		16'hB966: out_word = 8'hFE;
		16'hB967: out_word = 8'h80;
		16'hB968: out_word = 8'h20;
		16'hB969: out_word = 8'h05;
		16'hB96A: out_word = 8'h21;
		16'hB96B: out_word = 8'h0F;
		16'hB96C: out_word = 8'h27;
		16'hB96D: out_word = 8'h18;
		16'hB96E: out_word = 8'h11;
		16'hB96F: out_word = 8'h22;
		16'hB970: out_word = 8'h77;
		16'hB971: out_word = 8'h5B;
		16'hB972: out_word = 8'hCD;
		16'hB973: out_word = 8'h0B;
		16'hB974: out_word = 8'h3A;
		16'hB975: out_word = 8'h2A;
		16'hB976: out_word = 8'h96;
		16'hB977: out_word = 8'h5B;
		16'hB978: out_word = 8'hEF;
		16'hB979: out_word = 8'hA9;
		16'hB97A: out_word = 8'h30;
		16'hB97B: out_word = 8'hED;
		16'hB97C: out_word = 8'h5B;
		16'hB97D: out_word = 8'h94;
		16'hB97E: out_word = 8'h5B;
		16'hB97F: out_word = 8'h19;
		16'hB980: out_word = 8'h11;
		16'hB981: out_word = 8'h73;
		16'hB982: out_word = 8'h5B;
		16'hB983: out_word = 8'hE5;
		16'hB984: out_word = 8'hCD;
		16'hB985: out_word = 8'h3C;
		16'hB986: out_word = 8'h3A;
		16'hB987: out_word = 8'h58;
		16'hB988: out_word = 8'h1C;
		16'hB989: out_word = 8'h16;
		16'hB98A: out_word = 8'h00;
		16'hB98B: out_word = 8'hD5;
		16'hB98C: out_word = 8'hE5;
		16'hB98D: out_word = 8'h6B;
		16'hB98E: out_word = 8'h26;
		16'hB98F: out_word = 8'h00;
		16'hB990: out_word = 8'hED;
		16'hB991: out_word = 8'h4B;
		16'hB992: out_word = 8'h71;
		16'hB993: out_word = 8'h5B;
		16'hB994: out_word = 8'hB7;
		16'hB995: out_word = 8'hED;
		16'hB996: out_word = 8'h42;
		16'hB997: out_word = 8'h22;
		16'hB998: out_word = 8'h71;
		16'hB999: out_word = 8'h5B;
		16'hB99A: out_word = 8'h28;
		16'hB99B: out_word = 8'h33;
		16'hB99C: out_word = 8'h38;
		16'hB99D: out_word = 8'h27;
		16'hB99E: out_word = 8'h44;
		16'hB99F: out_word = 8'h4D;
		16'hB9A0: out_word = 8'h2A;
		16'hB9A1: out_word = 8'h79;
		16'hB9A2: out_word = 8'h5B;
		16'hB9A3: out_word = 8'hE5;
		16'hB9A4: out_word = 8'hD5;
		16'hB9A5: out_word = 8'h2A;
		16'hB9A6: out_word = 8'h65;
		16'hB9A7: out_word = 8'h5C;
		16'hB9A8: out_word = 8'h09;
		16'hB9A9: out_word = 8'h38;
		16'hB9AA: out_word = 8'h13;
		16'hB9AB: out_word = 8'hEB;
		16'hB9AC: out_word = 8'h21;
		16'hB9AD: out_word = 8'h82;
		16'hB9AE: out_word = 8'h00;
		16'hB9AF: out_word = 8'h19;
		16'hB9B0: out_word = 8'h38;
		16'hB9B1: out_word = 8'h0C;
		16'hB9B2: out_word = 8'hED;
		16'hB9B3: out_word = 8'h72;
		16'hB9B4: out_word = 8'h3F;
		16'hB9B5: out_word = 8'h38;
		16'hB9B6: out_word = 8'h07;
		16'hB9B7: out_word = 8'hD1;
		16'hB9B8: out_word = 8'hE1;
		16'hB9B9: out_word = 8'hEF;
		16'hB9BA: out_word = 8'h55;
		16'hB9BB: out_word = 8'h16;
		16'hB9BC: out_word = 8'h18;
		16'hB9BD: out_word = 8'h11;
		16'hB9BE: out_word = 8'hD1;
		16'hB9BF: out_word = 8'hE1;
		16'hB9C0: out_word = 8'hCD;
		16'hB9C1: out_word = 8'h45;
		16'hB9C2: out_word = 8'h1F;
		16'hB9C3: out_word = 8'hA7;
		16'hB9C4: out_word = 8'hC9;
		16'hB9C5: out_word = 8'h0B;
		16'hB9C6: out_word = 8'h1D;
		16'hB9C7: out_word = 8'h20;
		16'hB9C8: out_word = 8'hFC;
		16'hB9C9: out_word = 8'h2A;
		16'hB9CA: out_word = 8'h79;
		16'hB9CB: out_word = 8'h5B;
		16'hB9CC: out_word = 8'hEF;
		16'hB9CD: out_word = 8'hE8;
		16'hB9CE: out_word = 8'h19;
		16'hB9CF: out_word = 8'hED;
		16'hB9D0: out_word = 8'h5B;
		16'hB9D1: out_word = 8'h79;
		16'hB9D2: out_word = 8'h5B;
		16'hB9D3: out_word = 8'hE1;
		16'hB9D4: out_word = 8'hC1;
		16'hB9D5: out_word = 8'hED;
		16'hB9D6: out_word = 8'hB0;
		16'hB9D7: out_word = 8'hEB;
		16'hB9D8: out_word = 8'h36;
		16'hB9D9: out_word = 8'h0E;
		16'hB9DA: out_word = 8'hC1;
		16'hB9DB: out_word = 8'h23;
		16'hB9DC: out_word = 8'hE5;
		16'hB9DD: out_word = 8'hEF;
		16'hB9DE: out_word = 8'h2B;
		16'hB9DF: out_word = 8'h2D;
		16'hB9E0: out_word = 8'hD1;
		16'hB9E1: out_word = 8'h01;
		16'hB9E2: out_word = 8'h05;
		16'hB9E3: out_word = 8'h00;
		16'hB9E4: out_word = 8'hED;
		16'hB9E5: out_word = 8'hB0;
		16'hB9E6: out_word = 8'hEB;
		16'hB9E7: out_word = 8'hE5;
		16'hB9E8: out_word = 8'h2A;
		16'hB9E9: out_word = 8'h92;
		16'hB9EA: out_word = 8'h5B;
		16'hB9EB: out_word = 8'hE5;
		16'hB9EC: out_word = 8'h5E;
		16'hB9ED: out_word = 8'h23;
		16'hB9EE: out_word = 8'h56;
		16'hB9EF: out_word = 8'h2A;
		16'hB9F0: out_word = 8'h71;
		16'hB9F1: out_word = 8'h5B;
		16'hB9F2: out_word = 8'h19;
		16'hB9F3: out_word = 8'hEB;
		16'hB9F4: out_word = 8'hE1;
		16'hB9F5: out_word = 8'h73;
		16'hB9F6: out_word = 8'h23;
		16'hB9F7: out_word = 8'h72;
		16'hB9F8: out_word = 8'h2A;
		16'hB9F9: out_word = 8'h6B;
		16'hB9FA: out_word = 8'h5B;
		16'hB9FB: out_word = 8'hED;
		16'hB9FC: out_word = 8'h5B;
		16'hB9FD: out_word = 8'h71;
		16'hB9FE: out_word = 8'h5B;
		16'hB9FF: out_word = 8'h19;
		16'hBA00: out_word = 8'h22;
		16'hBA01: out_word = 8'h6B;
		16'hBA02: out_word = 8'h5B;
		16'hBA03: out_word = 8'hE1;
		16'hBA04: out_word = 8'hC9;
		16'hBA05: out_word = 8'h2A;
		16'hBA06: out_word = 8'h4B;
		16'hBA07: out_word = 8'h5C;
		16'hBA08: out_word = 8'h22;
		16'hBA09: out_word = 8'h77;
		16'hBA0A: out_word = 8'h5B;
		16'hBA0B: out_word = 8'h2A;
		16'hBA0C: out_word = 8'h53;
		16'hBA0D: out_word = 8'h5C;
		16'hBA0E: out_word = 8'hED;
		16'hBA0F: out_word = 8'h5B;
		16'hBA10: out_word = 8'h77;
		16'hBA11: out_word = 8'h5B;
		16'hBA12: out_word = 8'hB7;
		16'hBA13: out_word = 8'hED;
		16'hBA14: out_word = 8'h52;
		16'hBA15: out_word = 8'h28;
		16'hBA16: out_word = 8'h1A;
		16'hBA17: out_word = 8'h2A;
		16'hBA18: out_word = 8'h53;
		16'hBA19: out_word = 8'h5C;
		16'hBA1A: out_word = 8'h01;
		16'hBA1B: out_word = 8'h00;
		16'hBA1C: out_word = 8'h00;
		16'hBA1D: out_word = 8'hC5;
		16'hBA1E: out_word = 8'hEF;
		16'hBA1F: out_word = 8'hB8;
		16'hBA20: out_word = 8'h19;
		16'hBA21: out_word = 8'h2A;
		16'hBA22: out_word = 8'h77;
		16'hBA23: out_word = 8'h5B;
		16'hBA24: out_word = 8'hA7;
		16'hBA25: out_word = 8'hED;
		16'hBA26: out_word = 8'h52;
		16'hBA27: out_word = 8'h28;
		16'hBA28: out_word = 8'h05;
		16'hBA29: out_word = 8'hEB;
		16'hBA2A: out_word = 8'hC1;
		16'hBA2B: out_word = 8'h03;
		16'hBA2C: out_word = 8'h18;
		16'hBA2D: out_word = 8'hEF;
		16'hBA2E: out_word = 8'hD1;
		16'hBA2F: out_word = 8'h13;
		16'hBA30: out_word = 8'hC9;
		16'hBA31: out_word = 8'h11;
		16'hBA32: out_word = 8'h00;
		16'hBA33: out_word = 8'h00;
		16'hBA34: out_word = 8'hC9;
		16'hBA35: out_word = 8'h23;
		16'hBA36: out_word = 8'h7E;
		16'hBA37: out_word = 8'hFE;
		16'hBA38: out_word = 8'h20;
		16'hBA39: out_word = 8'h28;
		16'hBA3A: out_word = 8'hFA;
		16'hBA3B: out_word = 8'hC9;
		16'hBA3C: out_word = 8'hD5;
		16'hBA3D: out_word = 8'h01;
		16'hBA3E: out_word = 8'h18;
		16'hBA3F: out_word = 8'hFC;
		16'hBA40: out_word = 8'hCD;
		16'hBA41: out_word = 8'h60;
		16'hBA42: out_word = 8'h3A;
		16'hBA43: out_word = 8'h01;
		16'hBA44: out_word = 8'h9C;
		16'hBA45: out_word = 8'hFF;
		16'hBA46: out_word = 8'hCD;
		16'hBA47: out_word = 8'h60;
		16'hBA48: out_word = 8'h3A;
		16'hBA49: out_word = 8'h0E;
		16'hBA4A: out_word = 8'hF6;
		16'hBA4B: out_word = 8'hCD;
		16'hBA4C: out_word = 8'h60;
		16'hBA4D: out_word = 8'h3A;
		16'hBA4E: out_word = 8'h7D;
		16'hBA4F: out_word = 8'hC6;
		16'hBA50: out_word = 8'h30;
		16'hBA51: out_word = 8'h12;
		16'hBA52: out_word = 8'h13;
		16'hBA53: out_word = 8'h06;
		16'hBA54: out_word = 8'h03;
		16'hBA55: out_word = 8'hE1;
		16'hBA56: out_word = 8'h7E;
		16'hBA57: out_word = 8'hFE;
		16'hBA58: out_word = 8'h30;
		16'hBA59: out_word = 8'hC0;
		16'hBA5A: out_word = 8'h36;
		16'hBA5B: out_word = 8'h20;
		16'hBA5C: out_word = 8'h23;
		16'hBA5D: out_word = 8'h10;
		16'hBA5E: out_word = 8'hF7;
		16'hBA5F: out_word = 8'hC9;
		16'hBA60: out_word = 8'hAF;
		16'hBA61: out_word = 8'h09;
		16'hBA62: out_word = 8'h3C;
		16'hBA63: out_word = 8'h38;
		16'hBA64: out_word = 8'hFC;
		16'hBA65: out_word = 8'hED;
		16'hBA66: out_word = 8'h42;
		16'hBA67: out_word = 8'h3D;
		16'hBA68: out_word = 8'hC6;
		16'hBA69: out_word = 8'h30;
		16'hBA6A: out_word = 8'h12;
		16'hBA6B: out_word = 8'h13;
		16'hBA6C: out_word = 8'hC9;
		16'hBA6D: out_word = 8'h08;
		16'hBA6E: out_word = 8'h00;
		16'hBA6F: out_word = 8'h00;
		16'hBA70: out_word = 8'h14;
		16'hBA71: out_word = 8'h00;
		16'hBA72: out_word = 8'h00;
		16'hBA73: out_word = 8'h00;
		16'hBA74: out_word = 8'h0F;
		16'hBA75: out_word = 8'h00;
		16'hBA76: out_word = 8'h08;
		16'hBA77: out_word = 8'h00;
		16'hBA78: out_word = 8'h16;
		16'hBA79: out_word = 8'h01;
		16'hBA7A: out_word = 8'h00;
		16'hBA7B: out_word = 8'h00;
		16'hBA7C: out_word = 8'h00;
		16'hBA7D: out_word = 8'h0F;
		16'hBA7E: out_word = 8'h00;
		16'hBA7F: out_word = 8'hDD;
		16'hBA80: out_word = 8'h21;
		16'hBA81: out_word = 8'h6C;
		16'hBA82: out_word = 8'hFD;
		16'hBA83: out_word = 8'h21;
		16'hBA84: out_word = 8'h6D;
		16'hBA85: out_word = 8'h3A;
		16'hBA86: out_word = 8'h18;
		16'hBA87: out_word = 8'h03;
		16'hBA88: out_word = 8'h21;
		16'hBA89: out_word = 8'h76;
		16'hBA8A: out_word = 8'h3A;
		16'hBA8B: out_word = 8'h11;
		16'hBA8C: out_word = 8'h6C;
		16'hBA8D: out_word = 8'hFD;
		16'hBA8E: out_word = 8'hC3;
		16'hBA8F: out_word = 8'hBA;
		16'hBA90: out_word = 8'h3F;
		16'hBA91: out_word = 8'hD7;
		16'hBA92: out_word = 8'h7A;
		16'hBA93: out_word = 8'hD7;
		16'hBA94: out_word = 8'h37;
		16'hBA95: out_word = 8'hC9;
		16'hBA96: out_word = 8'hE6;
		16'hBA97: out_word = 8'h3F;
		16'hBA98: out_word = 8'hDD;
		16'hBA99: out_word = 8'h77;
		16'hBA9A: out_word = 8'h06;
		16'hBA9B: out_word = 8'h37;
		16'hBA9C: out_word = 8'hC9;
		16'hBA9D: out_word = 8'hDD;
		16'hBA9E: out_word = 8'h7E;
		16'hBA9F: out_word = 8'h01;
		16'hBAA0: out_word = 8'h80;
		16'hBAA1: out_word = 8'h47;
		16'hBAA2: out_word = 8'hCD;
		16'hBAA3: out_word = 8'hA0;
		16'hBAA4: out_word = 8'h3B;
		16'hBAA5: out_word = 8'h7E;
		16'hBAA6: out_word = 8'hDD;
		16'hBAA7: out_word = 8'h77;
		16'hBAA8: out_word = 8'h07;
		16'hBAA9: out_word = 8'h2F;
		16'hBAAA: out_word = 8'hE6;
		16'hBAAB: out_word = 8'hC0;
		16'hBAAC: out_word = 8'hDD;
		16'hBAAD: out_word = 8'hB6;
		16'hBAAE: out_word = 8'h06;
		16'hBAAF: out_word = 8'h77;
		16'hBAB0: out_word = 8'h37;
		16'hBAB1: out_word = 8'hC9;
		16'hBAB2: out_word = 8'hDD;
		16'hBAB3: out_word = 8'h7E;
		16'hBAB4: out_word = 8'h01;
		16'hBAB5: out_word = 8'h80;
		16'hBAB6: out_word = 8'h47;
		16'hBAB7: out_word = 8'hCD;
		16'hBAB8: out_word = 8'hA0;
		16'hBAB9: out_word = 8'h3B;
		16'hBABA: out_word = 8'hDD;
		16'hBABB: out_word = 8'h7E;
		16'hBABC: out_word = 8'h07;
		16'hBABD: out_word = 8'h77;
		16'hBABE: out_word = 8'hC9;
		16'hBABF: out_word = 8'hE5;
		16'hBAC0: out_word = 8'h26;
		16'hBAC1: out_word = 8'h00;
		16'hBAC2: out_word = 8'h7B;
		16'hBAC3: out_word = 8'h90;
		16'hBAC4: out_word = 8'h18;
		16'hBAC5: out_word = 8'h07;
		16'hBAC6: out_word = 8'hE5;
		16'hBAC7: out_word = 8'h7B;
		16'hBAC8: out_word = 8'h58;
		16'hBAC9: out_word = 8'h47;
		16'hBACA: out_word = 8'h93;
		16'hBACB: out_word = 8'h26;
		16'hBACC: out_word = 8'hFF;
		16'hBACD: out_word = 8'h4F;
		16'hBACE: out_word = 8'h78;
		16'hBACF: out_word = 8'hBB;
		16'hBAD0: out_word = 8'h28;
		16'hBAD1: out_word = 8'h4B;
		16'hBAD2: out_word = 8'hD5;
		16'hBAD3: out_word = 8'hCD;
		16'hBAD4: out_word = 8'h98;
		16'hBAD5: out_word = 8'h3B;
		16'hBAD6: out_word = 8'hC5;
		16'hBAD7: out_word = 8'h4C;
		16'hBAD8: out_word = 8'hEF;
		16'hBAD9: out_word = 8'h9B;
		16'hBADA: out_word = 8'h0E;
		16'hBADB: out_word = 8'hEB;
		16'hBADC: out_word = 8'hAF;
		16'hBADD: out_word = 8'hB1;
		16'hBADE: out_word = 8'h28;
		16'hBADF: out_word = 8'h03;
		16'hBAE0: out_word = 8'h04;
		16'hBAE1: out_word = 8'h18;
		16'hBAE2: out_word = 8'h01;
		16'hBAE3: out_word = 8'h05;
		16'hBAE4: out_word = 8'hD5;
		16'hBAE5: out_word = 8'hEF;
		16'hBAE6: out_word = 8'h9B;
		16'hBAE7: out_word = 8'h0E;
		16'hBAE8: out_word = 8'hD1;
		16'hBAE9: out_word = 8'h79;
		16'hBAEA: out_word = 8'h0E;
		16'hBAEB: out_word = 8'h20;
		16'hBAEC: out_word = 8'h06;
		16'hBAED: out_word = 8'h08;
		16'hBAEE: out_word = 8'hC5;
		16'hBAEF: out_word = 8'hE5;
		16'hBAF0: out_word = 8'hD5;
		16'hBAF1: out_word = 8'h06;
		16'hBAF2: out_word = 8'h00;
		16'hBAF3: out_word = 8'hED;
		16'hBAF4: out_word = 8'hB0;
		16'hBAF5: out_word = 8'hD1;
		16'hBAF6: out_word = 8'hE1;
		16'hBAF7: out_word = 8'hC1;
		16'hBAF8: out_word = 8'h24;
		16'hBAF9: out_word = 8'h14;
		16'hBAFA: out_word = 8'h10;
		16'hBAFB: out_word = 8'hF2;
		16'hBAFC: out_word = 8'hF5;
		16'hBAFD: out_word = 8'hD5;
		16'hBAFE: out_word = 8'hEF;
		16'hBAFF: out_word = 8'h88;
		16'hBB00: out_word = 8'h0E;
		16'hBB01: out_word = 8'hEB;
		16'hBB02: out_word = 8'hE3;
		16'hBB03: out_word = 8'hEF;
		16'hBB04: out_word = 8'h88;
		16'hBB05: out_word = 8'h0E;
		16'hBB06: out_word = 8'hEB;
		16'hBB07: out_word = 8'hE3;
		16'hBB08: out_word = 8'hD1;
		16'hBB09: out_word = 8'h01;
		16'hBB0A: out_word = 8'h20;
		16'hBB0B: out_word = 8'h00;
		16'hBB0C: out_word = 8'hED;
		16'hBB0D: out_word = 8'hB0;
		16'hBB0E: out_word = 8'hF1;
		16'hBB0F: out_word = 8'hC1;
		16'hBB10: out_word = 8'hA7;
		16'hBB11: out_word = 8'h28;
		16'hBB12: out_word = 8'h03;
		16'hBB13: out_word = 8'h04;
		16'hBB14: out_word = 8'h18;
		16'hBB15: out_word = 8'h01;
		16'hBB16: out_word = 8'h05;
		16'hBB17: out_word = 8'h0D;
		16'hBB18: out_word = 8'h67;
		16'hBB19: out_word = 8'h20;
		16'hBB1A: out_word = 8'hBB;
		16'hBB1B: out_word = 8'hD1;
		16'hBB1C: out_word = 8'h43;
		16'hBB1D: out_word = 8'hE1;
		16'hBB1E: out_word = 8'hCD;
		16'hBB1F: out_word = 8'hB8;
		16'hBB20: out_word = 8'h3B;
		16'hBB21: out_word = 8'hEB;
		16'hBB22: out_word = 8'h3A;
		16'hBB23: out_word = 8'h3C;
		16'hBB24: out_word = 8'h5C;
		16'hBB25: out_word = 8'hF5;
		16'hBB26: out_word = 8'h21;
		16'hBB27: out_word = 8'h0D;
		16'hBB28: out_word = 8'hEC;
		16'hBB29: out_word = 8'hCB;
		16'hBB2A: out_word = 8'h76;
		16'hBB2B: out_word = 8'hCB;
		16'hBB2C: out_word = 8'h87;
		16'hBB2D: out_word = 8'h28;
		16'hBB2E: out_word = 8'h02;
		16'hBB2F: out_word = 8'hCB;
		16'hBB30: out_word = 8'hC7;
		16'hBB31: out_word = 8'h32;
		16'hBB32: out_word = 8'h3C;
		16'hBB33: out_word = 8'h5C;
		16'hBB34: out_word = 8'h0E;
		16'hBB35: out_word = 8'h00;
		16'hBB36: out_word = 8'hCD;
		16'hBB37: out_word = 8'h2B;
		16'hBB38: out_word = 8'h37;
		16'hBB39: out_word = 8'hEB;
		16'hBB3A: out_word = 8'h06;
		16'hBB3B: out_word = 8'h20;
		16'hBB3C: out_word = 8'h7E;
		16'hBB3D: out_word = 8'hA7;
		16'hBB3E: out_word = 8'h20;
		16'hBB3F: out_word = 8'h02;
		16'hBB40: out_word = 8'h3E;
		16'hBB41: out_word = 8'h20;
		16'hBB42: out_word = 8'hFE;
		16'hBB43: out_word = 8'h90;
		16'hBB44: out_word = 8'h30;
		16'hBB45: out_word = 8'h0F;
		16'hBB46: out_word = 8'hEF;
		16'hBB47: out_word = 8'h10;
		16'hBB48: out_word = 8'h00;
		16'hBB49: out_word = 8'h23;
		16'hBB4A: out_word = 8'h10;
		16'hBB4B: out_word = 8'hF0;
		16'hBB4C: out_word = 8'hF1;
		16'hBB4D: out_word = 8'h32;
		16'hBB4E: out_word = 8'h3C;
		16'hBB4F: out_word = 8'h5C;
		16'hBB50: out_word = 8'hCD;
		16'hBB51: out_word = 8'hB8;
		16'hBB52: out_word = 8'h3B;
		16'hBB53: out_word = 8'h37;
		16'hBB54: out_word = 8'hC9;
		16'hBB55: out_word = 8'hCD;
		16'hBB56: out_word = 8'h20;
		16'hBB57: out_word = 8'h1F;
		16'hBB58: out_word = 8'hD7;
		16'hBB59: out_word = 8'hCD;
		16'hBB5A: out_word = 8'h45;
		16'hBB5B: out_word = 8'h1F;
		16'hBB5C: out_word = 8'h18;
		16'hBB5D: out_word = 8'hEB;
		16'hBB5E: out_word = 8'hCD;
		16'hBB5F: out_word = 8'hB8;
		16'hBB60: out_word = 8'h3B;
		16'hBB61: out_word = 8'h7A;
		16'hBB62: out_word = 8'h90;
		16'hBB63: out_word = 8'h3C;
		16'hBB64: out_word = 8'h4F;
		16'hBB65: out_word = 8'hCD;
		16'hBB66: out_word = 8'h98;
		16'hBB67: out_word = 8'h3B;
		16'hBB68: out_word = 8'hC5;
		16'hBB69: out_word = 8'hEF;
		16'hBB6A: out_word = 8'h9B;
		16'hBB6B: out_word = 8'h0E;
		16'hBB6C: out_word = 8'h0E;
		16'hBB6D: out_word = 8'h08;
		16'hBB6E: out_word = 8'hE5;
		16'hBB6F: out_word = 8'h06;
		16'hBB70: out_word = 8'h20;
		16'hBB71: out_word = 8'hAF;
		16'hBB72: out_word = 8'h77;
		16'hBB73: out_word = 8'h23;
		16'hBB74: out_word = 8'h10;
		16'hBB75: out_word = 8'hFC;
		16'hBB76: out_word = 8'hE1;
		16'hBB77: out_word = 8'h24;
		16'hBB78: out_word = 8'h0D;
		16'hBB79: out_word = 8'h20;
		16'hBB7A: out_word = 8'hF3;
		16'hBB7B: out_word = 8'h06;
		16'hBB7C: out_word = 8'h20;
		16'hBB7D: out_word = 8'hC5;
		16'hBB7E: out_word = 8'hEF;
		16'hBB7F: out_word = 8'h88;
		16'hBB80: out_word = 8'h0E;
		16'hBB81: out_word = 8'hEB;
		16'hBB82: out_word = 8'hC1;
		16'hBB83: out_word = 8'h3A;
		16'hBB84: out_word = 8'h8D;
		16'hBB85: out_word = 8'h5C;
		16'hBB86: out_word = 8'h77;
		16'hBB87: out_word = 8'h23;
		16'hBB88: out_word = 8'h10;
		16'hBB89: out_word = 8'hFC;
		16'hBB8A: out_word = 8'hC1;
		16'hBB8B: out_word = 8'h05;
		16'hBB8C: out_word = 8'h0D;
		16'hBB8D: out_word = 8'h20;
		16'hBB8E: out_word = 8'hD9;
		16'hBB8F: out_word = 8'hCD;
		16'hBB90: out_word = 8'hB8;
		16'hBB91: out_word = 8'h3B;
		16'hBB92: out_word = 8'h37;
		16'hBB93: out_word = 8'hC9;
		16'hBB94: out_word = 8'h3E;
		16'hBB95: out_word = 8'h21;
		16'hBB96: out_word = 8'h91;
		16'hBB97: out_word = 8'h4F;
		16'hBB98: out_word = 8'h3E;
		16'hBB99: out_word = 8'h18;
		16'hBB9A: out_word = 8'h90;
		16'hBB9B: out_word = 8'hDD;
		16'hBB9C: out_word = 8'h96;
		16'hBB9D: out_word = 8'h01;
		16'hBB9E: out_word = 8'h47;
		16'hBB9F: out_word = 8'hC9;
		16'hBBA0: out_word = 8'hC5;
		16'hBBA1: out_word = 8'hAF;
		16'hBBA2: out_word = 8'h50;
		16'hBBA3: out_word = 8'h5F;
		16'hBBA4: out_word = 8'hCB;
		16'hBBA5: out_word = 8'h1A;
		16'hBBA6: out_word = 8'hCB;
		16'hBBA7: out_word = 8'h1B;
		16'hBBA8: out_word = 8'hCB;
		16'hBBA9: out_word = 8'h1A;
		16'hBBAA: out_word = 8'hCB;
		16'hBBAB: out_word = 8'h1B;
		16'hBBAC: out_word = 8'hCB;
		16'hBBAD: out_word = 8'h1A;
		16'hBBAE: out_word = 8'hCB;
		16'hBBAF: out_word = 8'h1B;
		16'hBBB0: out_word = 8'h21;
		16'hBBB1: out_word = 8'h00;
		16'hBBB2: out_word = 8'h58;
		16'hBBB3: out_word = 8'h47;
		16'hBBB4: out_word = 8'h09;
		16'hBBB5: out_word = 8'h19;
		16'hBBB6: out_word = 8'hC1;
		16'hBBB7: out_word = 8'hC9;
		16'hBBB8: out_word = 8'hF5;
		16'hBBB9: out_word = 8'hE5;
		16'hBBBA: out_word = 8'hD5;
		16'hBBBB: out_word = 8'h2A;
		16'hBBBC: out_word = 8'h8D;
		16'hBBBD: out_word = 8'h5C;
		16'hBBBE: out_word = 8'hED;
		16'hBBBF: out_word = 8'h5B;
		16'hBBC0: out_word = 8'h8F;
		16'hBBC1: out_word = 8'h5C;
		16'hBBC2: out_word = 8'hD9;
		16'hBBC3: out_word = 8'h2A;
		16'hBBC4: out_word = 8'h0F;
		16'hBBC5: out_word = 8'hEC;
		16'hBBC6: out_word = 8'hED;
		16'hBBC7: out_word = 8'h5B;
		16'hBBC8: out_word = 8'h11;
		16'hBBC9: out_word = 8'hEC;
		16'hBBCA: out_word = 8'h22;
		16'hBBCB: out_word = 8'h8D;
		16'hBBCC: out_word = 8'h5C;
		16'hBBCD: out_word = 8'hED;
		16'hBBCE: out_word = 8'h53;
		16'hBBCF: out_word = 8'h8F;
		16'hBBD0: out_word = 8'h5C;
		16'hBBD1: out_word = 8'hD9;
		16'hBBD2: out_word = 8'h22;
		16'hBBD3: out_word = 8'h0F;
		16'hBBD4: out_word = 8'hEC;
		16'hBBD5: out_word = 8'hED;
		16'hBBD6: out_word = 8'h53;
		16'hBBD7: out_word = 8'h11;
		16'hBBD8: out_word = 8'hEC;
		16'hBBD9: out_word = 8'h21;
		16'hBBDA: out_word = 8'h13;
		16'hBBDB: out_word = 8'hEC;
		16'hBBDC: out_word = 8'h3A;
		16'hBBDD: out_word = 8'h91;
		16'hBBDE: out_word = 8'h5C;
		16'hBBDF: out_word = 8'h56;
		16'hBBE0: out_word = 8'h77;
		16'hBBE1: out_word = 8'h7A;
		16'hBBE2: out_word = 8'h32;
		16'hBBE3: out_word = 8'h91;
		16'hBBE4: out_word = 8'h5C;
		16'hBBE5: out_word = 8'hD1;
		16'hBBE6: out_word = 8'hE1;
		16'hBBE7: out_word = 8'hF1;
		16'hBBE8: out_word = 8'hC9;
		16'hBBE9: out_word = 8'hCD;
		16'hBBEA: out_word = 8'h56;
		16'hBBEB: out_word = 8'h3C;
		16'hBBEC: out_word = 8'h21;
		16'hBBED: out_word = 8'h3C;
		16'hBBEE: out_word = 8'h5C;
		16'hBBEF: out_word = 8'hCB;
		16'hBBF0: out_word = 8'h86;
		16'hBBF1: out_word = 8'hCB;
		16'hBBF2: out_word = 8'hF6;
		16'hBBF3: out_word = 8'h21;
		16'hBBF4: out_word = 8'h0E;
		16'hBBF5: out_word = 8'hEC;
		16'hBBF6: out_word = 8'h36;
		16'hBBF7: out_word = 8'hFF;
		16'hBBF8: out_word = 8'hCD;
		16'hBBF9: out_word = 8'h20;
		16'hBBFA: out_word = 8'h1F;
		16'hBBFB: out_word = 8'hEF;
		16'hBBFC: out_word = 8'hB0;
		16'hBBFD: out_word = 8'h16;
		16'hBBFE: out_word = 8'h2A;
		16'hBBFF: out_word = 8'h59;
		16'hBC00: out_word = 8'h5C;
		16'hBC01: out_word = 8'h01;
		16'hBC02: out_word = 8'h0A;
		16'hBC03: out_word = 8'h00;
		16'hBC04: out_word = 8'hEF;
		16'hBC05: out_word = 8'h55;
		16'hBC06: out_word = 8'h16;
		16'hBC07: out_word = 8'h21;
		16'hBC08: out_word = 8'h16;
		16'hBC09: out_word = 8'h3C;
		16'hBC0A: out_word = 8'hED;
		16'hBC0B: out_word = 8'h5B;
		16'hBC0C: out_word = 8'h59;
		16'hBC0D: out_word = 8'h5C;
		16'hBC0E: out_word = 8'h01;
		16'hBC0F: out_word = 8'h0A;
		16'hBC10: out_word = 8'h00;
		16'hBC11: out_word = 8'hED;
		16'hBC12: out_word = 8'hB0;
		16'hBC13: out_word = 8'hC3;
		16'hBC14: out_word = 8'h11;
		16'hBC15: out_word = 8'h1B;
		16'hBC16: out_word = 8'hF9;
		16'hBC17: out_word = 8'hC0;
		16'hBC18: out_word = 8'hB0;
		16'hBC19: out_word = 8'h22;
		16'hBC1A: out_word = 8'h31;
		16'hBC1B: out_word = 8'h35;
		16'hBC1C: out_word = 8'h36;
		16'hBC1D: out_word = 8'h31;
		16'hBC1E: out_word = 8'h36;
		16'hBC1F: out_word = 8'h22;
		16'hBC20: out_word = 8'h28;
		16'hBC21: out_word = 8'h09;
		16'hBC22: out_word = 8'hDB;
		16'hBC23: out_word = 8'hFE;
		16'hBC24: out_word = 8'hE6;
		16'hBC25: out_word = 8'h40;
		16'hBC26: out_word = 8'h28;
		16'hBC27: out_word = 8'hF5;
		16'hBC28: out_word = 8'h23;
		16'hBC29: out_word = 8'h18;
		16'hBC2A: out_word = 8'hF2;
		16'hBC2B: out_word = 8'hCB;
		16'hBC2C: out_word = 8'h15;
		16'hBC2D: out_word = 8'hCB;
		16'hBC2E: out_word = 8'h14;
		16'hBC2F: out_word = 8'hCB;
		16'hBC30: out_word = 8'h15;
		16'hBC31: out_word = 8'hCB;
		16'hBC32: out_word = 8'h14;
		16'hBC33: out_word = 8'h08;
		16'hBC34: out_word = 8'h28;
		16'hBC35: out_word = 8'h07;
		16'hBC36: out_word = 8'h08;
		16'hBC37: out_word = 8'h3E;
		16'hBC38: out_word = 8'h20;
		16'hBC39: out_word = 8'h94;
		16'hBC3A: out_word = 8'h6F;
		16'hBC3B: out_word = 8'h18;
		16'hBC3C: out_word = 8'h02;
		16'hBC3D: out_word = 8'h08;
		16'hBC3E: out_word = 8'h6C;
		16'hBC3F: out_word = 8'hAF;
		16'hBC40: out_word = 8'h67;
		16'hBC41: out_word = 8'h11;
		16'hBC42: out_word = 8'h1F;
		16'hBC43: out_word = 8'h59;
		16'hBC44: out_word = 8'h06;
		16'hBC45: out_word = 8'h20;
		16'hBC46: out_word = 8'h3E;
		16'hBC47: out_word = 8'h48;
		16'hBC48: out_word = 8'hFB;
		16'hBC49: out_word = 8'h76;
		16'hBC4A: out_word = 8'hF3;
		16'hBC4B: out_word = 8'h12;
		16'hBC4C: out_word = 8'h1B;
		16'hBC4D: out_word = 8'h10;
		16'hBC4E: out_word = 8'hFC;
		16'hBC4F: out_word = 8'h13;
		16'hBC50: out_word = 8'h19;
		16'hBC51: out_word = 8'h3E;
		16'hBC52: out_word = 8'h68;
		16'hBC53: out_word = 8'h77;
		16'hBC54: out_word = 8'h18;
		16'hBC55: out_word = 8'hA8;
		16'hBC56: out_word = 8'hFB;
		16'hBC57: out_word = 8'h06;
		16'hBC58: out_word = 8'h19;
		16'hBC59: out_word = 8'h76;
		16'hBC5A: out_word = 8'h10;
		16'hBC5B: out_word = 8'hFD;
		16'hBC5C: out_word = 8'h21;
		16'hBC5D: out_word = 8'h3B;
		16'hBC5E: out_word = 8'h5C;
		16'hBC5F: out_word = 8'hCB;
		16'hBC60: out_word = 8'hAE;
		16'hBC61: out_word = 8'h37;
		16'hBC62: out_word = 8'hC9;
		16'hBC63: out_word = 8'h3E;
		16'hBC64: out_word = 8'h01;
		16'hBC65: out_word = 8'h18;
		16'hBC66: out_word = 8'h02;
		16'hBC67: out_word = 8'h3E;
		16'hBC68: out_word = 8'h00;
		16'hBC69: out_word = 8'h32;
		16'hBC6A: out_word = 8'h8A;
		16'hBC6B: out_word = 8'hFD;
		16'hBC6C: out_word = 8'h21;
		16'hBC6D: out_word = 8'h00;
		16'hBC6E: out_word = 8'h00;
		16'hBC6F: out_word = 8'h22;
		16'hBC70: out_word = 8'h85;
		16'hBC71: out_word = 8'hFD;
		16'hBC72: out_word = 8'h22;
		16'hBC73: out_word = 8'h87;
		16'hBC74: out_word = 8'hFD;
		16'hBC75: out_word = 8'h39;
		16'hBC76: out_word = 8'h22;
		16'hBC77: out_word = 8'h8B;
		16'hBC78: out_word = 8'hFD;
		16'hBC79: out_word = 8'hCD;
		16'hBC7A: out_word = 8'hEA;
		16'hBC7B: out_word = 8'h34;
		16'hBC7C: out_word = 8'h3E;
		16'hBC7D: out_word = 8'h00;
		16'hBC7E: out_word = 8'h32;
		16'hBC7F: out_word = 8'h84;
		16'hBC80: out_word = 8'hFD;
		16'hBC81: out_word = 8'h21;
		16'hBC82: out_word = 8'h74;
		16'hBC83: out_word = 8'hFD;
		16'hBC84: out_word = 8'h22;
		16'hBC85: out_word = 8'h7D;
		16'hBC86: out_word = 8'hFD;
		16'hBC87: out_word = 8'hCD;
		16'hBC88: out_word = 8'h20;
		16'hBC89: out_word = 8'h1F;
		16'hBC8A: out_word = 8'hEF;
		16'hBC8B: out_word = 8'hB0;
		16'hBC8C: out_word = 8'h16;
		16'hBC8D: out_word = 8'hCD;
		16'hBC8E: out_word = 8'h45;
		16'hBC8F: out_word = 8'h1F;
		16'hBC90: out_word = 8'h3E;
		16'hBC91: out_word = 8'h00;
		16'hBC92: out_word = 8'h32;
		16'hBC93: out_word = 8'h81;
		16'hBC94: out_word = 8'hFD;
		16'hBC95: out_word = 8'h2A;
		16'hBC96: out_word = 8'h59;
		16'hBC97: out_word = 8'h5C;
		16'hBC98: out_word = 8'h22;
		16'hBC99: out_word = 8'h82;
		16'hBC9A: out_word = 8'hFD;
		16'hBC9B: out_word = 8'h21;
		16'hBC9C: out_word = 8'h00;
		16'hBC9D: out_word = 8'h00;
		16'hBC9E: out_word = 8'h22;
		16'hBC9F: out_word = 8'h7F;
		16'hBCA0: out_word = 8'hFD;
		16'hBCA1: out_word = 8'h2A;
		16'hBCA2: out_word = 8'h85;
		16'hBCA3: out_word = 8'hFD;
		16'hBCA4: out_word = 8'h23;
		16'hBCA5: out_word = 8'h22;
		16'hBCA6: out_word = 8'h85;
		16'hBCA7: out_word = 8'hFD;
		16'hBCA8: out_word = 8'hCD;
		16'hBCA9: out_word = 8'h9D;
		16'hBCAA: out_word = 8'h3D;
		16'hBCAB: out_word = 8'h4F;
		16'hBCAC: out_word = 8'h3A;
		16'hBCAD: out_word = 8'h81;
		16'hBCAE: out_word = 8'hFD;
		16'hBCAF: out_word = 8'hFE;
		16'hBCB0: out_word = 8'h00;
		16'hBCB1: out_word = 8'h20;
		16'hBCB2: out_word = 8'h41;
		16'hBCB3: out_word = 8'h79;
		16'hBCB4: out_word = 8'hE6;
		16'hBCB5: out_word = 8'h04;
		16'hBCB6: out_word = 8'h28;
		16'hBCB7: out_word = 8'h35;
		16'hBCB8: out_word = 8'hCD;
		16'hBCB9: out_word = 8'hE9;
		16'hBCBA: out_word = 8'h3D;
		16'hBCBB: out_word = 8'h30;
		16'hBCBC: out_word = 8'h07;
		16'hBCBD: out_word = 8'h3E;
		16'hBCBE: out_word = 8'h01;
		16'hBCBF: out_word = 8'h32;
		16'hBCC0: out_word = 8'h81;
		16'hBCC1: out_word = 8'hFD;
		16'hBCC2: out_word = 8'h18;
		16'hBCC3: out_word = 8'hDD;
		16'hBCC4: out_word = 8'h2A;
		16'hBCC5: out_word = 8'h7F;
		16'hBCC6: out_word = 8'hFD;
		16'hBCC7: out_word = 8'h7D;
		16'hBCC8: out_word = 8'hB4;
		16'hBCC9: out_word = 8'hC2;
		16'hBCCA: out_word = 8'h1E;
		16'hBCCB: out_word = 8'h3D;
		16'hBCCC: out_word = 8'hC5;
		16'hBCCD: out_word = 8'hCD;
		16'hBCCE: out_word = 8'hCD;
		16'hBCCF: out_word = 8'h3D;
		16'hBCD0: out_word = 8'hC1;
		16'hBCD1: out_word = 8'h3E;
		16'hBCD2: out_word = 8'h00;
		16'hBCD3: out_word = 8'h32;
		16'hBCD4: out_word = 8'h81;
		16'hBCD5: out_word = 8'hFD;
		16'hBCD6: out_word = 8'h79;
		16'hBCD7: out_word = 8'hE6;
		16'hBCD8: out_word = 8'h01;
		16'hBCD9: out_word = 8'h20;
		16'hBCDA: out_word = 8'hD8;
		16'hBCDB: out_word = 8'h78;
		16'hBCDC: out_word = 8'hCD;
		16'hBCDD: out_word = 8'h16;
		16'hBCDE: out_word = 8'h3E;
		16'hBCDF: out_word = 8'hD0;
		16'hBCE0: out_word = 8'h2A;
		16'hBCE1: out_word = 8'h85;
		16'hBCE2: out_word = 8'hFD;
		16'hBCE3: out_word = 8'h23;
		16'hBCE4: out_word = 8'h22;
		16'hBCE5: out_word = 8'h85;
		16'hBCE6: out_word = 8'hFD;
		16'hBCE7: out_word = 8'hCD;
		16'hBCE8: out_word = 8'h9D;
		16'hBCE9: out_word = 8'h3D;
		16'hBCEA: out_word = 8'h4F;
		16'hBCEB: out_word = 8'h18;
		16'hBCEC: out_word = 8'hE9;
		16'hBCED: out_word = 8'h78;
		16'hBCEE: out_word = 8'hCD;
		16'hBCEF: out_word = 8'h16;
		16'hBCF0: out_word = 8'h3E;
		16'hBCF1: out_word = 8'hD0;
		16'hBCF2: out_word = 8'h18;
		16'hBCF3: out_word = 8'hAD;
		16'hBCF4: out_word = 8'hFE;
		16'hBCF5: out_word = 8'h01;
		16'hBCF6: out_word = 8'h20;
		16'hBCF7: out_word = 8'hF5;
		16'hBCF8: out_word = 8'h79;
		16'hBCF9: out_word = 8'hE6;
		16'hBCFA: out_word = 8'h01;
		16'hBCFB: out_word = 8'h28;
		16'hBCFC: out_word = 8'hBB;
		16'hBCFD: out_word = 8'hC5;
		16'hBCFE: out_word = 8'hCD;
		16'hBCFF: out_word = 8'h7E;
		16'hBD00: out_word = 8'h3F;
		16'hBD01: out_word = 8'hC1;
		16'hBD02: out_word = 8'h38;
		16'hBD03: out_word = 8'h79;
		16'hBD04: out_word = 8'h2A;
		16'hBD05: out_word = 8'h7F;
		16'hBD06: out_word = 8'hFD;
		16'hBD07: out_word = 8'h7C;
		16'hBD08: out_word = 8'hB5;
		16'hBD09: out_word = 8'h20;
		16'hBD0A: out_word = 8'h13;
		16'hBD0B: out_word = 8'h79;
		16'hBD0C: out_word = 8'hE6;
		16'hBD0D: out_word = 8'h02;
		16'hBD0E: out_word = 8'h28;
		16'hBD0F: out_word = 8'hBC;
		16'hBD10: out_word = 8'hCD;
		16'hBD11: out_word = 8'hE9;
		16'hBD12: out_word = 8'h3D;
		16'hBD13: out_word = 8'h30;
		16'hBD14: out_word = 8'hAF;
		16'hBD15: out_word = 8'h2A;
		16'hBD16: out_word = 8'h7D;
		16'hBD17: out_word = 8'hFD;
		16'hBD18: out_word = 8'h2B;
		16'hBD19: out_word = 8'h22;
		16'hBD1A: out_word = 8'h7F;
		16'hBD1B: out_word = 8'hFD;
		16'hBD1C: out_word = 8'h18;
		16'hBD1D: out_word = 8'h83;
		16'hBD1E: out_word = 8'hC5;
		16'hBD1F: out_word = 8'h21;
		16'hBD20: out_word = 8'h74;
		16'hBD21: out_word = 8'hFD;
		16'hBD22: out_word = 8'hED;
		16'hBD23: out_word = 8'h5B;
		16'hBD24: out_word = 8'h7F;
		16'hBD25: out_word = 8'hFD;
		16'hBD26: out_word = 8'h7A;
		16'hBD27: out_word = 8'hBC;
		16'hBD28: out_word = 8'h20;
		16'hBD29: out_word = 8'h05;
		16'hBD2A: out_word = 8'h7B;
		16'hBD2B: out_word = 8'hBD;
		16'hBD2C: out_word = 8'h20;
		16'hBD2D: out_word = 8'h01;
		16'hBD2E: out_word = 8'h13;
		16'hBD2F: out_word = 8'h1B;
		16'hBD30: out_word = 8'h18;
		16'hBD31: out_word = 8'h01;
		16'hBD32: out_word = 8'h23;
		16'hBD33: out_word = 8'h7E;
		16'hBD34: out_word = 8'hE6;
		16'hBD35: out_word = 8'h7F;
		16'hBD36: out_word = 8'hE5;
		16'hBD37: out_word = 8'hD5;
		16'hBD38: out_word = 8'hCD;
		16'hBD39: out_word = 8'h16;
		16'hBD3A: out_word = 8'h3E;
		16'hBD3B: out_word = 8'hD1;
		16'hBD3C: out_word = 8'hE1;
		16'hBD3D: out_word = 8'h7C;
		16'hBD3E: out_word = 8'hBA;
		16'hBD3F: out_word = 8'h20;
		16'hBD40: out_word = 8'hF1;
		16'hBD41: out_word = 8'h7D;
		16'hBD42: out_word = 8'hBB;
		16'hBD43: out_word = 8'h20;
		16'hBD44: out_word = 8'hED;
		16'hBD45: out_word = 8'hED;
		16'hBD46: out_word = 8'h5B;
		16'hBD47: out_word = 8'h7F;
		16'hBD48: out_word = 8'hFD;
		16'hBD49: out_word = 8'h21;
		16'hBD4A: out_word = 8'h74;
		16'hBD4B: out_word = 8'hFD;
		16'hBD4C: out_word = 8'h22;
		16'hBD4D: out_word = 8'h7F;
		16'hBD4E: out_word = 8'hFD;
		16'hBD4F: out_word = 8'hED;
		16'hBD50: out_word = 8'h4B;
		16'hBD51: out_word = 8'h7D;
		16'hBD52: out_word = 8'hFD;
		16'hBD53: out_word = 8'h0B;
		16'hBD54: out_word = 8'h7A;
		16'hBD55: out_word = 8'hBC;
		16'hBD56: out_word = 8'h20;
		16'hBD57: out_word = 8'h18;
		16'hBD58: out_word = 8'h7B;
		16'hBD59: out_word = 8'hBD;
		16'hBD5A: out_word = 8'h20;
		16'hBD5B: out_word = 8'h14;
		16'hBD5C: out_word = 8'h13;
		16'hBD5D: out_word = 8'hE5;
		16'hBD5E: out_word = 8'h21;
		16'hBD5F: out_word = 8'h00;
		16'hBD60: out_word = 8'h00;
		16'hBD61: out_word = 8'h22;
		16'hBD62: out_word = 8'h7F;
		16'hBD63: out_word = 8'hFD;
		16'hBD64: out_word = 8'hE1;
		16'hBD65: out_word = 8'h78;
		16'hBD66: out_word = 8'hBC;
		16'hBD67: out_word = 8'h20;
		16'hBD68: out_word = 8'h07;
		16'hBD69: out_word = 8'h79;
		16'hBD6A: out_word = 8'hBD;
		16'hBD6B: out_word = 8'h20;
		16'hBD6C: out_word = 8'h03;
		16'hBD6D: out_word = 8'hC1;
		16'hBD6E: out_word = 8'h18;
		16'hBD6F: out_word = 8'h1F;
		16'hBD70: out_word = 8'h1A;
		16'hBD71: out_word = 8'h77;
		16'hBD72: out_word = 8'h23;
		16'hBD73: out_word = 8'h13;
		16'hBD74: out_word = 8'hE6;
		16'hBD75: out_word = 8'h80;
		16'hBD76: out_word = 8'h28;
		16'hBD77: out_word = 8'hF8;
		16'hBD78: out_word = 8'h22;
		16'hBD79: out_word = 8'h7D;
		16'hBD7A: out_word = 8'hFD;
		16'hBD7B: out_word = 8'h18;
		16'hBD7C: out_word = 8'h81;
		16'hBD7D: out_word = 8'hC5;
		16'hBD7E: out_word = 8'hCD;
		16'hBD7F: out_word = 8'h16;
		16'hBD80: out_word = 8'h3E;
		16'hBD81: out_word = 8'hC1;
		16'hBD82: out_word = 8'h21;
		16'hBD83: out_word = 8'h00;
		16'hBD84: out_word = 8'h00;
		16'hBD85: out_word = 8'h22;
		16'hBD86: out_word = 8'h7F;
		16'hBD87: out_word = 8'hFD;
		16'hBD88: out_word = 8'h3A;
		16'hBD89: out_word = 8'h81;
		16'hBD8A: out_word = 8'hFD;
		16'hBD8B: out_word = 8'hFE;
		16'hBD8C: out_word = 8'h04;
		16'hBD8D: out_word = 8'h28;
		16'hBD8E: out_word = 8'h05;
		16'hBD8F: out_word = 8'h3E;
		16'hBD90: out_word = 8'h00;
		16'hBD91: out_word = 8'h32;
		16'hBD92: out_word = 8'h81;
		16'hBD93: out_word = 8'hFD;
		16'hBD94: out_word = 8'h21;
		16'hBD95: out_word = 8'h74;
		16'hBD96: out_word = 8'hFD;
		16'hBD97: out_word = 8'h22;
		16'hBD98: out_word = 8'h7D;
		16'hBD99: out_word = 8'hFD;
		16'hBD9A: out_word = 8'hC3;
		16'hBD9B: out_word = 8'hB3;
		16'hBD9C: out_word = 8'h3C;
		16'hBD9D: out_word = 8'hCD;
		16'hBD9E: out_word = 8'h54;
		16'hBD9F: out_word = 8'h2D;
		16'hBDA0: out_word = 8'h47;
		16'hBDA1: out_word = 8'hFE;
		16'hBDA2: out_word = 8'h3F;
		16'hBDA3: out_word = 8'h38;
		16'hBDA4: out_word = 8'h0A;
		16'hBDA5: out_word = 8'hF6;
		16'hBDA6: out_word = 8'h20;
		16'hBDA7: out_word = 8'hCD;
		16'hBDA8: out_word = 8'hC6;
		16'hBDA9: out_word = 8'h3D;
		16'hBDAA: out_word = 8'h38;
		16'hBDAB: out_word = 8'h17;
		16'hBDAC: out_word = 8'h3E;
		16'hBDAD: out_word = 8'h01;
		16'hBDAE: out_word = 8'hC9;
		16'hBDAF: out_word = 8'hFE;
		16'hBDB0: out_word = 8'h20;
		16'hBDB1: out_word = 8'h28;
		16'hBDB2: out_word = 8'h0D;
		16'hBDB3: out_word = 8'hFE;
		16'hBDB4: out_word = 8'h23;
		16'hBDB5: out_word = 8'h28;
		16'hBDB6: out_word = 8'h06;
		16'hBDB7: out_word = 8'h38;
		16'hBDB8: out_word = 8'hF3;
		16'hBDB9: out_word = 8'hFE;
		16'hBDBA: out_word = 8'h24;
		16'hBDBB: out_word = 8'h20;
		16'hBDBC: out_word = 8'hEF;
		16'hBDBD: out_word = 8'h3E;
		16'hBDBE: out_word = 8'h02;
		16'hBDBF: out_word = 8'hC9;
		16'hBDC0: out_word = 8'h3E;
		16'hBDC1: out_word = 8'h03;
		16'hBDC2: out_word = 8'hC9;
		16'hBDC3: out_word = 8'h3E;
		16'hBDC4: out_word = 8'h06;
		16'hBDC5: out_word = 8'hC9;
		16'hBDC6: out_word = 8'hFE;
		16'hBDC7: out_word = 8'h7B;
		16'hBDC8: out_word = 8'hD0;
		16'hBDC9: out_word = 8'hFE;
		16'hBDCA: out_word = 8'h61;
		16'hBDCB: out_word = 8'h3F;
		16'hBDCC: out_word = 8'hC9;
		16'hBDCD: out_word = 8'h21;
		16'hBDCE: out_word = 8'h74;
		16'hBDCF: out_word = 8'hFD;
		16'hBDD0: out_word = 8'h22;
		16'hBDD1: out_word = 8'h7D;
		16'hBDD2: out_word = 8'hFD;
		16'hBDD3: out_word = 8'h97;
		16'hBDD4: out_word = 8'h32;
		16'hBDD5: out_word = 8'h7F;
		16'hBDD6: out_word = 8'hFD;
		16'hBDD7: out_word = 8'h32;
		16'hBDD8: out_word = 8'h80;
		16'hBDD9: out_word = 8'hFD;
		16'hBDDA: out_word = 8'h7E;
		16'hBDDB: out_word = 8'hE6;
		16'hBDDC: out_word = 8'h7F;
		16'hBDDD: out_word = 8'hE5;
		16'hBDDE: out_word = 8'hCD;
		16'hBDDF: out_word = 8'h9C;
		16'hBDE0: out_word = 8'h3E;
		16'hBDE1: out_word = 8'hE1;
		16'hBDE2: out_word = 8'h7E;
		16'hBDE3: out_word = 8'hE6;
		16'hBDE4: out_word = 8'h80;
		16'hBDE5: out_word = 8'hC0;
		16'hBDE6: out_word = 8'h23;
		16'hBDE7: out_word = 8'h18;
		16'hBDE8: out_word = 8'hF1;
		16'hBDE9: out_word = 8'h2A;
		16'hBDEA: out_word = 8'h7D;
		16'hBDEB: out_word = 8'hFD;
		16'hBDEC: out_word = 8'h11;
		16'hBDED: out_word = 8'h7D;
		16'hBDEE: out_word = 8'hFD;
		16'hBDEF: out_word = 8'h7A;
		16'hBDF0: out_word = 8'hBC;
		16'hBDF1: out_word = 8'h20;
		16'hBDF2: out_word = 8'h05;
		16'hBDF3: out_word = 8'h7B;
		16'hBDF4: out_word = 8'hBD;
		16'hBDF5: out_word = 8'hCA;
		16'hBDF6: out_word = 8'h13;
		16'hBDF7: out_word = 8'h3E;
		16'hBDF8: out_word = 8'h11;
		16'hBDF9: out_word = 8'h74;
		16'hBDFA: out_word = 8'hFD;
		16'hBDFB: out_word = 8'h7A;
		16'hBDFC: out_word = 8'hBC;
		16'hBDFD: out_word = 8'h20;
		16'hBDFE: out_word = 8'h04;
		16'hBDFF: out_word = 8'h7B;
		16'hBE00: out_word = 8'hBD;
		16'hBE01: out_word = 8'h28;
		16'hBE02: out_word = 8'h06;
		16'hBE03: out_word = 8'h2B;
		16'hBE04: out_word = 8'h7E;
		16'hBE05: out_word = 8'hE6;
		16'hBE06: out_word = 8'h7F;
		16'hBE07: out_word = 8'h77;
		16'hBE08: out_word = 8'h23;
		16'hBE09: out_word = 8'h78;
		16'hBE0A: out_word = 8'hF6;
		16'hBE0B: out_word = 8'h80;
		16'hBE0C: out_word = 8'h77;
		16'hBE0D: out_word = 8'h23;
		16'hBE0E: out_word = 8'h22;
		16'hBE0F: out_word = 8'h7D;
		16'hBE10: out_word = 8'hFD;
		16'hBE11: out_word = 8'h37;
		16'hBE12: out_word = 8'hC9;
		16'hBE13: out_word = 8'h37;
		16'hBE14: out_word = 8'h3F;
		16'hBE15: out_word = 8'hC9;
		16'hBE16: out_word = 8'hF5;
		16'hBE17: out_word = 8'h3A;
		16'hBE18: out_word = 8'h89;
		16'hBE19: out_word = 8'hFD;
		16'hBE1A: out_word = 8'hB7;
		16'hBE1B: out_word = 8'h20;
		16'hBE1C: out_word = 8'h12;
		16'hBE1D: out_word = 8'hF1;
		16'hBE1E: out_word = 8'hFE;
		16'hBE1F: out_word = 8'h3E;
		16'hBE20: out_word = 8'h28;
		16'hBE21: out_word = 8'h08;
		16'hBE22: out_word = 8'hFE;
		16'hBE23: out_word = 8'h3C;
		16'hBE24: out_word = 8'h28;
		16'hBE25: out_word = 8'h04;
		16'hBE26: out_word = 8'hCD;
		16'hBE27: out_word = 8'h64;
		16'hBE28: out_word = 8'h3E;
		16'hBE29: out_word = 8'hC9;
		16'hBE2A: out_word = 8'h32;
		16'hBE2B: out_word = 8'h89;
		16'hBE2C: out_word = 8'hFD;
		16'hBE2D: out_word = 8'h37;
		16'hBE2E: out_word = 8'hC9;
		16'hBE2F: out_word = 8'hFE;
		16'hBE30: out_word = 8'h3C;
		16'hBE31: out_word = 8'h3E;
		16'hBE32: out_word = 8'h00;
		16'hBE33: out_word = 8'h32;
		16'hBE34: out_word = 8'h89;
		16'hBE35: out_word = 8'hFD;
		16'hBE36: out_word = 8'h20;
		16'hBE37: out_word = 8'h1A;
		16'hBE38: out_word = 8'hF1;
		16'hBE39: out_word = 8'hFE;
		16'hBE3A: out_word = 8'h3E;
		16'hBE3B: out_word = 8'h20;
		16'hBE3C: out_word = 8'h04;
		16'hBE3D: out_word = 8'h3E;
		16'hBE3E: out_word = 8'hC9;
		16'hBE3F: out_word = 8'h18;
		16'hBE40: out_word = 8'hE5;
		16'hBE41: out_word = 8'hFE;
		16'hBE42: out_word = 8'h3D;
		16'hBE43: out_word = 8'h20;
		16'hBE44: out_word = 8'h04;
		16'hBE45: out_word = 8'h3E;
		16'hBE46: out_word = 8'hC7;
		16'hBE47: out_word = 8'h18;
		16'hBE48: out_word = 8'hDD;
		16'hBE49: out_word = 8'hF5;
		16'hBE4A: out_word = 8'h3E;
		16'hBE4B: out_word = 8'h3C;
		16'hBE4C: out_word = 8'hCD;
		16'hBE4D: out_word = 8'h64;
		16'hBE4E: out_word = 8'h3E;
		16'hBE4F: out_word = 8'hF1;
		16'hBE50: out_word = 8'h18;
		16'hBE51: out_word = 8'hD4;
		16'hBE52: out_word = 8'hF1;
		16'hBE53: out_word = 8'hFE;
		16'hBE54: out_word = 8'h3D;
		16'hBE55: out_word = 8'h20;
		16'hBE56: out_word = 8'h04;
		16'hBE57: out_word = 8'h3E;
		16'hBE58: out_word = 8'hC8;
		16'hBE59: out_word = 8'h18;
		16'hBE5A: out_word = 8'hCB;
		16'hBE5B: out_word = 8'hF5;
		16'hBE5C: out_word = 8'h3E;
		16'hBE5D: out_word = 8'h3E;
		16'hBE5E: out_word = 8'hCD;
		16'hBE5F: out_word = 8'h64;
		16'hBE60: out_word = 8'h3E;
		16'hBE61: out_word = 8'hF1;
		16'hBE62: out_word = 8'h18;
		16'hBE63: out_word = 8'hC2;
		16'hBE64: out_word = 8'hFE;
		16'hBE65: out_word = 8'h0D;
		16'hBE66: out_word = 8'h28;
		16'hBE67: out_word = 8'h20;
		16'hBE68: out_word = 8'hFE;
		16'hBE69: out_word = 8'hEA;
		16'hBE6A: out_word = 8'h47;
		16'hBE6B: out_word = 8'h20;
		16'hBE6C: out_word = 8'h07;
		16'hBE6D: out_word = 8'h3E;
		16'hBE6E: out_word = 8'h04;
		16'hBE6F: out_word = 8'h32;
		16'hBE70: out_word = 8'h81;
		16'hBE71: out_word = 8'hFD;
		16'hBE72: out_word = 8'h18;
		16'hBE73: out_word = 8'h0E;
		16'hBE74: out_word = 8'hFE;
		16'hBE75: out_word = 8'h22;
		16'hBE76: out_word = 8'h20;
		16'hBE77: out_word = 8'h0A;
		16'hBE78: out_word = 8'h3A;
		16'hBE79: out_word = 8'h81;
		16'hBE7A: out_word = 8'hFD;
		16'hBE7B: out_word = 8'hE6;
		16'hBE7C: out_word = 8'hFE;
		16'hBE7D: out_word = 8'hEE;
		16'hBE7E: out_word = 8'h02;
		16'hBE7F: out_word = 8'h32;
		16'hBE80: out_word = 8'h81;
		16'hBE81: out_word = 8'hFD;
		16'hBE82: out_word = 8'h78;
		16'hBE83: out_word = 8'hCD;
		16'hBE84: out_word = 8'h9C;
		16'hBE85: out_word = 8'h3E;
		16'hBE86: out_word = 8'h37;
		16'hBE87: out_word = 8'hC9;
		16'hBE88: out_word = 8'h3A;
		16'hBE89: out_word = 8'h8A;
		16'hBE8A: out_word = 8'hFD;
		16'hBE8B: out_word = 8'hFE;
		16'hBE8C: out_word = 8'h00;
		16'hBE8D: out_word = 8'h28;
		16'hBE8E: out_word = 8'h0A;
		16'hBE8F: out_word = 8'hED;
		16'hBE90: out_word = 8'h4B;
		16'hBE91: out_word = 8'h85;
		16'hBE92: out_word = 8'hFD;
		16'hBE93: out_word = 8'h2A;
		16'hBE94: out_word = 8'h8B;
		16'hBE95: out_word = 8'hFD;
		16'hBE96: out_word = 8'hF9;
		16'hBE97: out_word = 8'h37;
		16'hBE98: out_word = 8'hC9;
		16'hBE99: out_word = 8'h37;
		16'hBE9A: out_word = 8'h3F;
		16'hBE9B: out_word = 8'hC9;
		16'hBE9C: out_word = 8'h5F;
		16'hBE9D: out_word = 8'h3A;
		16'hBE9E: out_word = 8'h84;
		16'hBE9F: out_word = 8'hFD;
		16'hBEA0: out_word = 8'h57;
		16'hBEA1: out_word = 8'h7B;
		16'hBEA2: out_word = 8'hFE;
		16'hBEA3: out_word = 8'h20;
		16'hBEA4: out_word = 8'h20;
		16'hBEA5: out_word = 8'h20;
		16'hBEA6: out_word = 8'h7A;
		16'hBEA7: out_word = 8'hE6;
		16'hBEA8: out_word = 8'h01;
		16'hBEA9: out_word = 8'h20;
		16'hBEAA: out_word = 8'h14;
		16'hBEAB: out_word = 8'h7A;
		16'hBEAC: out_word = 8'hE6;
		16'hBEAD: out_word = 8'h02;
		16'hBEAE: out_word = 8'h20;
		16'hBEAF: out_word = 8'h07;
		16'hBEB0: out_word = 8'h7A;
		16'hBEB1: out_word = 8'hF6;
		16'hBEB2: out_word = 8'h02;
		16'hBEB3: out_word = 8'h32;
		16'hBEB4: out_word = 8'h84;
		16'hBEB5: out_word = 8'hFD;
		16'hBEB6: out_word = 8'hC9;
		16'hBEB7: out_word = 8'h7B;
		16'hBEB8: out_word = 8'hCD;
		16'hBEB9: out_word = 8'hFB;
		16'hBEBA: out_word = 8'h3E;
		16'hBEBB: out_word = 8'h3A;
		16'hBEBC: out_word = 8'h84;
		16'hBEBD: out_word = 8'hFD;
		16'hBEBE: out_word = 8'hC9;
		16'hBEBF: out_word = 8'h7A;
		16'hBEC0: out_word = 8'hE6;
		16'hBEC1: out_word = 8'hFE;
		16'hBEC2: out_word = 8'h32;
		16'hBEC3: out_word = 8'h84;
		16'hBEC4: out_word = 8'hFD;
		16'hBEC5: out_word = 8'hC9;
		16'hBEC6: out_word = 8'hFE;
		16'hBEC7: out_word = 8'hA3;
		16'hBEC8: out_word = 8'h30;
		16'hBEC9: out_word = 8'h24;
		16'hBECA: out_word = 8'h7A;
		16'hBECB: out_word = 8'hE6;
		16'hBECC: out_word = 8'h02;
		16'hBECD: out_word = 8'h20;
		16'hBECE: out_word = 8'h0B;
		16'hBECF: out_word = 8'h7A;
		16'hBED0: out_word = 8'hE6;
		16'hBED1: out_word = 8'hFE;
		16'hBED2: out_word = 8'h32;
		16'hBED3: out_word = 8'h84;
		16'hBED4: out_word = 8'hFD;
		16'hBED5: out_word = 8'h7B;
		16'hBED6: out_word = 8'hCD;
		16'hBED7: out_word = 8'hFB;
		16'hBED8: out_word = 8'h3E;
		16'hBED9: out_word = 8'hC9;
		16'hBEDA: out_word = 8'hD5;
		16'hBEDB: out_word = 8'h3E;
		16'hBEDC: out_word = 8'h20;
		16'hBEDD: out_word = 8'hCD;
		16'hBEDE: out_word = 8'hFB;
		16'hBEDF: out_word = 8'h3E;
		16'hBEE0: out_word = 8'hD1;
		16'hBEE1: out_word = 8'h7A;
		16'hBEE2: out_word = 8'hE6;
		16'hBEE3: out_word = 8'hFE;
		16'hBEE4: out_word = 8'hE6;
		16'hBEE5: out_word = 8'hFD;
		16'hBEE6: out_word = 8'h32;
		16'hBEE7: out_word = 8'h84;
		16'hBEE8: out_word = 8'hFD;
		16'hBEE9: out_word = 8'h7B;
		16'hBEEA: out_word = 8'hCD;
		16'hBEEB: out_word = 8'hFB;
		16'hBEEC: out_word = 8'h3E;
		16'hBEED: out_word = 8'hC9;
		16'hBEEE: out_word = 8'h7A;
		16'hBEEF: out_word = 8'hE6;
		16'hBEF0: out_word = 8'hFD;
		16'hBEF1: out_word = 8'hF6;
		16'hBEF2: out_word = 8'h01;
		16'hBEF3: out_word = 8'h32;
		16'hBEF4: out_word = 8'h84;
		16'hBEF5: out_word = 8'hFD;
		16'hBEF6: out_word = 8'h7B;
		16'hBEF7: out_word = 8'hCD;
		16'hBEF8: out_word = 8'hFB;
		16'hBEF9: out_word = 8'h3E;
		16'hBEFA: out_word = 8'hC9;
		16'hBEFB: out_word = 8'h2A;
		16'hBEFC: out_word = 8'h87;
		16'hBEFD: out_word = 8'hFD;
		16'hBEFE: out_word = 8'h23;
		16'hBEFF: out_word = 8'h22;
		16'hBF00: out_word = 8'h87;
		16'hBF01: out_word = 8'hFD;
		16'hBF02: out_word = 8'h2A;
		16'hBF03: out_word = 8'h82;
		16'hBF04: out_word = 8'hFD;
		16'hBF05: out_word = 8'h47;
		16'hBF06: out_word = 8'h3A;
		16'hBF07: out_word = 8'h8A;
		16'hBF08: out_word = 8'hFD;
		16'hBF09: out_word = 8'hFE;
		16'hBF0A: out_word = 8'h00;
		16'hBF0B: out_word = 8'h78;
		16'hBF0C: out_word = 8'h28;
		16'hBF0D: out_word = 8'h25;
		16'hBF0E: out_word = 8'hED;
		16'hBF0F: out_word = 8'h5B;
		16'hBF10: out_word = 8'h5F;
		16'hBF11: out_word = 8'h5C;
		16'hBF12: out_word = 8'h7C;
		16'hBF13: out_word = 8'hBA;
		16'hBF14: out_word = 8'h20;
		16'hBF15: out_word = 8'h1A;
		16'hBF16: out_word = 8'h7D;
		16'hBF17: out_word = 8'hBB;
		16'hBF18: out_word = 8'h20;
		16'hBF19: out_word = 8'h16;
		16'hBF1A: out_word = 8'hED;
		16'hBF1B: out_word = 8'h4B;
		16'hBF1C: out_word = 8'h85;
		16'hBF1D: out_word = 8'hFD;
		16'hBF1E: out_word = 8'h2A;
		16'hBF1F: out_word = 8'h87;
		16'hBF20: out_word = 8'hFD;
		16'hBF21: out_word = 8'hA7;
		16'hBF22: out_word = 8'hED;
		16'hBF23: out_word = 8'h42;
		16'hBF24: out_word = 8'h30;
		16'hBF25: out_word = 8'h04;
		16'hBF26: out_word = 8'hED;
		16'hBF27: out_word = 8'h4B;
		16'hBF28: out_word = 8'h87;
		16'hBF29: out_word = 8'hFD;
		16'hBF2A: out_word = 8'h2A;
		16'hBF2B: out_word = 8'h8B;
		16'hBF2C: out_word = 8'hFD;
		16'hBF2D: out_word = 8'hF9;
		16'hBF2E: out_word = 8'h37;
		16'hBF2F: out_word = 8'hC9;
		16'hBF30: out_word = 8'h37;
		16'hBF31: out_word = 8'h18;
		16'hBF32: out_word = 8'h02;
		16'hBF33: out_word = 8'h37;
		16'hBF34: out_word = 8'h3F;
		16'hBF35: out_word = 8'hCD;
		16'hBF36: out_word = 8'h20;
		16'hBF37: out_word = 8'h1F;
		16'hBF38: out_word = 8'h30;
		16'hBF39: out_word = 8'h0D;
		16'hBF3A: out_word = 8'h7E;
		16'hBF3B: out_word = 8'hEB;
		16'hBF3C: out_word = 8'hFE;
		16'hBF3D: out_word = 8'h0E;
		16'hBF3E: out_word = 8'h20;
		16'hBF3F: out_word = 8'h1D;
		16'hBF40: out_word = 8'h13;
		16'hBF41: out_word = 8'h13;
		16'hBF42: out_word = 8'h13;
		16'hBF43: out_word = 8'h13;
		16'hBF44: out_word = 8'h13;
		16'hBF45: out_word = 8'h18;
		16'hBF46: out_word = 8'h16;
		16'hBF47: out_word = 8'hF5;
		16'hBF48: out_word = 8'h01;
		16'hBF49: out_word = 8'h01;
		16'hBF4A: out_word = 8'h00;
		16'hBF4B: out_word = 8'hE5;
		16'hBF4C: out_word = 8'hD5;
		16'hBF4D: out_word = 8'hCD;
		16'hBF4E: out_word = 8'h66;
		16'hBF4F: out_word = 8'h3F;
		16'hBF50: out_word = 8'hD1;
		16'hBF51: out_word = 8'hE1;
		16'hBF52: out_word = 8'hEF;
		16'hBF53: out_word = 8'h64;
		16'hBF54: out_word = 8'h16;
		16'hBF55: out_word = 8'h2A;
		16'hBF56: out_word = 8'h65;
		16'hBF57: out_word = 8'h5C;
		16'hBF58: out_word = 8'hEB;
		16'hBF59: out_word = 8'hED;
		16'hBF5A: out_word = 8'hB8;
		16'hBF5B: out_word = 8'hF1;
		16'hBF5C: out_word = 8'h12;
		16'hBF5D: out_word = 8'h13;
		16'hBF5E: out_word = 8'hCD;
		16'hBF5F: out_word = 8'h45;
		16'hBF60: out_word = 8'h1F;
		16'hBF61: out_word = 8'hED;
		16'hBF62: out_word = 8'h53;
		16'hBF63: out_word = 8'h82;
		16'hBF64: out_word = 8'hFD;
		16'hBF65: out_word = 8'hC9;
		16'hBF66: out_word = 8'h2A;
		16'hBF67: out_word = 8'h65;
		16'hBF68: out_word = 8'h5C;
		16'hBF69: out_word = 8'h09;
		16'hBF6A: out_word = 8'h38;
		16'hBF6B: out_word = 8'h0A;
		16'hBF6C: out_word = 8'hEB;
		16'hBF6D: out_word = 8'h21;
		16'hBF6E: out_word = 8'h82;
		16'hBF6F: out_word = 8'h00;
		16'hBF70: out_word = 8'h19;
		16'hBF71: out_word = 8'h38;
		16'hBF72: out_word = 8'h03;
		16'hBF73: out_word = 8'hED;
		16'hBF74: out_word = 8'h72;
		16'hBF75: out_word = 8'hD8;
		16'hBF76: out_word = 8'h3E;
		16'hBF77: out_word = 8'h03;
		16'hBF78: out_word = 8'h32;
		16'hBF79: out_word = 8'h3A;
		16'hBF7A: out_word = 8'h5C;
		16'hBF7B: out_word = 8'hC3;
		16'hBF7C: out_word = 8'h21;
		16'hBF7D: out_word = 8'h03;
		16'hBF7E: out_word = 8'hCD;
		16'hBF7F: out_word = 8'h2E;
		16'hBF80: out_word = 8'hFD;
		16'hBF81: out_word = 8'hD8;
		16'hBF82: out_word = 8'h06;
		16'hBF83: out_word = 8'hF9;
		16'hBF84: out_word = 8'h11;
		16'hBF85: out_word = 8'h74;
		16'hBF86: out_word = 8'hFD;
		16'hBF87: out_word = 8'h21;
		16'hBF88: out_word = 8'h94;
		16'hBF89: out_word = 8'h35;
		16'hBF8A: out_word = 8'hCD;
		16'hBF8B: out_word = 8'h3B;
		16'hBF8C: out_word = 8'hFD;
		16'hBF8D: out_word = 8'hD0;
		16'hBF8E: out_word = 8'hFE;
		16'hBF8F: out_word = 8'hFF;
		16'hBF90: out_word = 8'h20;
		16'hBF91: out_word = 8'h04;
		16'hBF92: out_word = 8'h3E;
		16'hBF93: out_word = 8'hD4;
		16'hBF94: out_word = 8'h18;
		16'hBF95: out_word = 8'h22;
		16'hBF96: out_word = 8'hFE;
		16'hBF97: out_word = 8'hFE;
		16'hBF98: out_word = 8'h20;
		16'hBF99: out_word = 8'h04;
		16'hBF9A: out_word = 8'h3E;
		16'hBF9B: out_word = 8'hD3;
		16'hBF9C: out_word = 8'h18;
		16'hBF9D: out_word = 8'h1A;
		16'hBF9E: out_word = 8'hFE;
		16'hBF9F: out_word = 8'hFD;
		16'hBFA0: out_word = 8'h20;
		16'hBFA1: out_word = 8'h04;
		16'hBFA2: out_word = 8'h3E;
		16'hBFA3: out_word = 8'hCE;
		16'hBFA4: out_word = 8'h18;
		16'hBFA5: out_word = 8'h12;
		16'hBFA6: out_word = 8'hFE;
		16'hBFA7: out_word = 8'hFC;
		16'hBFA8: out_word = 8'h20;
		16'hBFA9: out_word = 8'h04;
		16'hBFAA: out_word = 8'h3E;
		16'hBFAB: out_word = 8'hED;
		16'hBFAC: out_word = 8'h18;
		16'hBFAD: out_word = 8'h0A;
		16'hBFAE: out_word = 8'hFE;
		16'hBFAF: out_word = 8'hFB;
		16'hBFB0: out_word = 8'h20;
		16'hBFB1: out_word = 8'h04;
		16'hBFB2: out_word = 8'h3E;
		16'hBFB3: out_word = 8'hEC;
		16'hBFB4: out_word = 8'h18;
		16'hBFB5: out_word = 8'h02;
		16'hBFB6: out_word = 8'hD6;
		16'hBFB7: out_word = 8'h56;
		16'hBFB8: out_word = 8'h37;
		16'hBFB9: out_word = 8'hC9;
		16'hBFBA: out_word = 8'h46;
		16'hBFBB: out_word = 8'h23;
		16'hBFBC: out_word = 8'h7E;
		16'hBFBD: out_word = 8'h12;
		16'hBFBE: out_word = 8'h13;
		16'hBFBF: out_word = 8'h23;
		16'hBFC0: out_word = 8'h10;
		16'hBFC1: out_word = 8'hFA;
		16'hBFC2: out_word = 8'hC9;
		16'hBFC3: out_word = 8'hFE;
		16'hBFC4: out_word = 8'h30;
		16'hBFC5: out_word = 8'h3F;
		16'hBFC6: out_word = 8'hD0;
		16'hBFC7: out_word = 8'hFE;
		16'hBFC8: out_word = 8'h3A;
		16'hBFC9: out_word = 8'hD0;
		16'hBFCA: out_word = 8'hD6;
		16'hBFCB: out_word = 8'h30;
		16'hBFCC: out_word = 8'h37;
		16'hBFCD: out_word = 8'hC9;
		16'hBFCE: out_word = 8'hC5;
		16'hBFCF: out_word = 8'hD5;
		16'hBFD0: out_word = 8'h46;
		16'hBFD1: out_word = 8'h23;
		16'hBFD2: out_word = 8'hBE;
		16'hBFD3: out_word = 8'h23;
		16'hBFD4: out_word = 8'h5E;
		16'hBFD5: out_word = 8'h23;
		16'hBFD6: out_word = 8'h56;
		16'hBFD7: out_word = 8'h28;
		16'hBFD8: out_word = 8'h08;
		16'hBFD9: out_word = 8'h23;
		16'hBFDA: out_word = 8'h10;
		16'hBFDB: out_word = 8'hF6;
		16'hBFDC: out_word = 8'h37;
		16'hBFDD: out_word = 8'h3F;
		16'hBFDE: out_word = 8'hD1;
		16'hBFDF: out_word = 8'hC1;
		16'hBFE0: out_word = 8'hC9;
		16'hBFE1: out_word = 8'hEB;
		16'hBFE2: out_word = 8'hD1;
		16'hBFE3: out_word = 8'hC1;
		16'hBFE4: out_word = 8'hCD;
		16'hBFE5: out_word = 8'hEE;
		16'hBFE6: out_word = 8'h3F;
		16'hBFE7: out_word = 8'h38;
		16'hBFE8: out_word = 8'h02;
		16'hBFE9: out_word = 8'hBF;
		16'hBFEA: out_word = 8'hC9;
		16'hBFEB: out_word = 8'hBF;
		16'hBFEC: out_word = 8'h37;
		16'hBFED: out_word = 8'hC9;
		16'hBFEE: out_word = 8'hE9;
		16'hBFEF: out_word = 8'h00;
		16'hBFF0: out_word = 8'h4D;
		16'hBFF1: out_word = 8'h42;
		16'hBFF2: out_word = 8'h00;
		16'hBFF3: out_word = 8'h53;
		16'hBFF4: out_word = 8'h42;
		16'hBFF5: out_word = 8'h00;
		16'hBFF6: out_word = 8'h41;
		16'hBFF7: out_word = 8'h43;
		16'hBFF8: out_word = 8'h00;
		16'hBFF9: out_word = 8'h52;
		16'hBFFA: out_word = 8'h47;
		16'hBFFB: out_word = 8'h00;
		16'hBFFC: out_word = 8'h4B;
		16'hBFFD: out_word = 8'h4D;
		16'hBFFE: out_word = 8'h00;
		16'hBFFF: out_word = 8'h01;
		16'hC000: out_word = 8'hF3;
		16'hC001: out_word = 8'h31;
		16'hC002: out_word = 8'h00;
		16'hC003: out_word = 8'h60;
		16'hC004: out_word = 8'hFD;
		16'hC005: out_word = 8'h21;
		16'hC006: out_word = 8'h3A;
		16'hC007: out_word = 8'h5C;
		16'hC008: out_word = 8'h3E;
		16'hC009: out_word = 8'h3F;
		16'hC00A: out_word = 8'hED;
		16'hC00B: out_word = 8'h47;
		16'hC00C: out_word = 8'hED;
		16'hC00D: out_word = 8'h56;
		16'hC00E: out_word = 8'hAF;
		16'hC00F: out_word = 8'hD3;
		16'hC010: out_word = 8'hFE;
		16'hC011: out_word = 8'hDD;
		16'hC012: out_word = 8'h2E;
		16'hC013: out_word = 8'h50;
		16'hC014: out_word = 8'h21;
		16'hC015: out_word = 8'h04;
		16'hC016: out_word = 8'h00;
		16'hC017: out_word = 8'h16;
		16'hC018: out_word = 8'h40;
		16'hC019: out_word = 8'h5D;
		16'hC01A: out_word = 8'h06;
		16'hC01B: out_word = 8'h80;
		16'hC01C: out_word = 8'h4D;
		16'hC01D: out_word = 8'h0A;
		16'hC01E: out_word = 8'hBE;
		16'hC01F: out_word = 8'hC2;
		16'hC020: out_word = 8'h7D;
		16'hC021: out_word = 8'h00;
		16'hC022: out_word = 8'hEB;
		16'hC023: out_word = 8'hBE;
		16'hC024: out_word = 8'hEB;
		16'hC025: out_word = 8'hC2;
		16'hC026: out_word = 8'h7D;
		16'hC027: out_word = 8'h00;
		16'hC028: out_word = 8'h2D;
		16'hC029: out_word = 8'h1D;
		16'hC02A: out_word = 8'h0D;
		16'hC02B: out_word = 8'h20;
		16'hC02C: out_word = 8'hF0;
		16'hC02D: out_word = 8'hDD;
		16'hC02E: out_word = 8'h2E;
		16'hC02F: out_word = 8'h41;
		16'hC030: out_word = 8'h11;
		16'hC031: out_word = 8'h02;
		16'hC032: out_word = 8'h10;
		16'hC033: out_word = 8'h01;
		16'hC034: out_word = 8'h77;
		16'hC035: out_word = 8'h00;
		16'hC036: out_word = 8'hED;
		16'hC037: out_word = 8'h59;
		16'hC038: out_word = 8'h21;
		16'hC039: out_word = 8'hA6;
		16'hC03A: out_word = 8'h3F;
		16'hC03B: out_word = 8'h01;
		16'hC03C: out_word = 8'hFD;
		16'hC03D: out_word = 8'h7F;
		16'hC03E: out_word = 8'hED;
		16'hC03F: out_word = 8'h51;
		16'hC040: out_word = 8'h01;
		16'hC041: out_word = 8'hF7;
		16'hC042: out_word = 8'h3F;
		16'hC043: out_word = 8'h7E;
		16'hC044: out_word = 8'hED;
		16'hC045: out_word = 8'h79;
		16'hC046: out_word = 8'h23;
		16'hC047: out_word = 8'h78;
		16'hC048: out_word = 8'hC6;
		16'hC049: out_word = 8'h40;
		16'hC04A: out_word = 8'h47;
		16'hC04B: out_word = 8'h30;
		16'hC04C: out_word = 8'hF6;
		16'hC04D: out_word = 8'h7A;
		16'hC04E: out_word = 8'hEE;
		16'hC04F: out_word = 8'h10;
		16'hC050: out_word = 8'h57;
		16'hC051: out_word = 8'h28;
		16'hC052: out_word = 8'hE8;
		16'hC053: out_word = 8'h3E;
		16'hC054: out_word = 8'hAB;
		16'hC055: out_word = 8'h01;
		16'hC056: out_word = 8'h77;
		16'hC057: out_word = 8'h41;
		16'hC058: out_word = 8'hED;
		16'hC059: out_word = 8'h79;
		16'hC05A: out_word = 8'h21;
		16'hC05B: out_word = 8'hBE;
		16'hC05C: out_word = 8'h3F;
		16'hC05D: out_word = 8'h11;
		16'hC05E: out_word = 8'h0F;
		16'hC05F: out_word = 8'hAB;
		16'hC060: out_word = 8'h01;
		16'hC061: out_word = 8'h77;
		16'hC062: out_word = 8'h01;
		16'hC063: out_word = 8'hED;
		16'hC064: out_word = 8'h51;
		16'hC065: out_word = 8'h7B;
		16'hC066: out_word = 8'hCB;
		16'hC067: out_word = 8'h5B;
		16'hC068: out_word = 8'hD3;
		16'hC069: out_word = 8'hFE;
		16'hC06A: out_word = 8'h28;
		16'hC06B: out_word = 8'h02;
		16'hC06C: out_word = 8'hD3;
		16'hC06D: out_word = 8'hF6;
		16'hC06E: out_word = 8'h7E;
		16'hC06F: out_word = 8'h23;
		16'hC070: out_word = 8'hD3;
		16'hC071: out_word = 8'hFF;
		16'hC072: out_word = 8'h1D;
		16'hC073: out_word = 8'hF2;
		16'hC074: out_word = 8'h65;
		16'hC075: out_word = 8'h00;
		16'hC076: out_word = 8'h3E;
		16'hC077: out_word = 8'hAB;
		16'hC078: out_word = 8'h01;
		16'hC079: out_word = 8'h77;
		16'hC07A: out_word = 8'h41;
		16'hC07B: out_word = 8'hED;
		16'hC07C: out_word = 8'h79;
		16'hC07D: out_word = 8'h01;
		16'hC07E: out_word = 8'hFF;
		16'hC07F: out_word = 8'hFE;
		16'hC080: out_word = 8'h78;
		16'hC081: out_word = 8'hDB;
		16'hC082: out_word = 8'hFE;
		16'hC083: out_word = 8'h1F;
		16'hC084: out_word = 8'h38;
		16'hC085: out_word = 8'h01;
		16'hC086: out_word = 8'h0C;
		16'hC087: out_word = 8'h1F;
		16'hC088: out_word = 8'h38;
		16'hC089: out_word = 8'h01;
		16'hC08A: out_word = 8'h0C;
		16'hC08B: out_word = 8'h1F;
		16'hC08C: out_word = 8'h38;
		16'hC08D: out_word = 8'h01;
		16'hC08E: out_word = 8'h0C;
		16'hC08F: out_word = 8'h1F;
		16'hC090: out_word = 8'h38;
		16'hC091: out_word = 8'h01;
		16'hC092: out_word = 8'h0C;
		16'hC093: out_word = 8'h1F;
		16'hC094: out_word = 8'h38;
		16'hC095: out_word = 8'h01;
		16'hC096: out_word = 8'h0C;
		16'hC097: out_word = 8'hCB;
		16'hC098: out_word = 8'h00;
		16'hC099: out_word = 8'h38;
		16'hC09A: out_word = 8'hE5;
		16'hC09B: out_word = 8'h0D;
		16'hC09C: out_word = 8'hF2;
		16'hC09D: out_word = 8'hF6;
		16'hC09E: out_word = 8'h00;
		16'hC09F: out_word = 8'h11;
		16'hC0A0: out_word = 8'h00;
		16'hC0A1: out_word = 8'h00;
		16'hC0A2: out_word = 8'h01;
		16'hC0A3: out_word = 8'hFD;
		16'hC0A4: out_word = 8'h7F;
		16'hC0A5: out_word = 8'hD5;
		16'hC0A6: out_word = 8'h3E;
		16'hC0A7: out_word = 8'hFE;
		16'hC0A8: out_word = 8'hDB;
		16'hC0A9: out_word = 8'hFE;
		16'hC0AA: out_word = 8'h1F;
		16'hC0AB: out_word = 8'h3E;
		16'hC0AC: out_word = 8'h00;
		16'hC0AD: out_word = 8'hD2;
		16'hC0AE: out_word = 8'h14;
		16'hC0AF: out_word = 8'h01;
		16'hC0B0: out_word = 8'h3E;
		16'hC0B1: out_word = 8'h7F;
		16'hC0B2: out_word = 8'hDB;
		16'hC0B3: out_word = 8'hFE;
		16'hC0B4: out_word = 8'h57;
		16'hC0B5: out_word = 8'h1F;
		16'hC0B6: out_word = 8'h1F;
		16'hC0B7: out_word = 8'h3E;
		16'hC0B8: out_word = 8'h10;
		16'hC0B9: out_word = 8'hD2;
		16'hC0BA: out_word = 8'h14;
		16'hC0BB: out_word = 8'h01;
		16'hC0BC: out_word = 8'h7A;
		16'hC0BD: out_word = 8'h1F;
		16'hC0BE: out_word = 8'h38;
		16'hC0BF: out_word = 8'h09;
		16'hC0C0: out_word = 8'h3E;
		16'hC0C1: out_word = 8'h10;
		16'hC0C2: out_word = 8'h11;
		16'hC0C3: out_word = 8'h2F;
		16'hC0C4: out_word = 8'h3D;
		16'hC0C5: out_word = 8'hD5;
		16'hC0C6: out_word = 8'hC3;
		16'hC0C7: out_word = 8'h14;
		16'hC0C8: out_word = 8'h01;
		16'hC0C9: out_word = 8'h3E;
		16'hC0CA: out_word = 8'hFD;
		16'hC0CB: out_word = 8'hDB;
		16'hC0CC: out_word = 8'hFE;
		16'hC0CD: out_word = 8'hE6;
		16'hC0CE: out_word = 8'h04;
		16'hC0CF: out_word = 8'hCA;
		16'hC0D0: out_word = 8'h07;
		16'hC0D1: out_word = 8'h01;
		16'hC0D2: out_word = 8'h21;
		16'hC0D3: out_word = 8'h00;
		16'hC0D4: out_word = 8'h60;
		16'hC0D5: out_word = 8'hF9;
		16'hC0D6: out_word = 8'hEB;
		16'hC0D7: out_word = 8'h21;
		16'hC0D8: out_word = 8'hA7;
		16'hC0D9: out_word = 8'h07;
		16'hC0DA: out_word = 8'hCD;
		16'hC0DB: out_word = 8'h38;
		16'hC0DC: out_word = 8'h3F;
		16'hC0DD: out_word = 8'h21;
		16'hC0DE: out_word = 8'hBA;
		16'hC0DF: out_word = 8'h30;
		16'hC0E0: out_word = 8'h11;
		16'hC0E1: out_word = 8'h00;
		16'hC0E2: out_word = 8'hF8;
		16'hC0E3: out_word = 8'hCD;
		16'hC0E4: out_word = 8'h38;
		16'hC0E5: out_word = 8'h3F;
		16'hC0E6: out_word = 8'hAF;
		16'hC0E7: out_word = 8'hDB;
		16'hC0E8: out_word = 8'hFE;
		16'hC0E9: out_word = 8'h2F;
		16'hC0EA: out_word = 8'hE6;
		16'hC0EB: out_word = 8'h1F;
		16'hC0EC: out_word = 8'h3E;
		16'hC0ED: out_word = 8'h10;
		16'hC0EE: out_word = 8'h20;
		16'hC0EF: out_word = 8'h09;
		16'hC0F0: out_word = 8'h21;
		16'hC0F1: out_word = 8'h00;
		16'hC0F2: out_word = 8'h60;
		16'hC0F3: out_word = 8'hE5;
		16'hC0F4: out_word = 8'h18;
		16'hC0F5: out_word = 8'h1E;
		16'hC0F6: out_word = 8'h37;
		16'hC0F7: out_word = 8'h3E;
		16'hC0F8: out_word = 8'h10;
		16'hC0F9: out_word = 8'h21;
		16'hC0FA: out_word = 8'h48;
		16'hC0FB: out_word = 8'h01;
		16'hC0FC: out_word = 8'h11;
		16'hC0FD: out_word = 8'h00;
		16'hC0FE: out_word = 8'h60;
		16'hC0FF: out_word = 8'hD5;
		16'hC100: out_word = 8'hF5;
		16'hC101: out_word = 8'hCD;
		16'hC102: out_word = 8'h38;
		16'hC103: out_word = 8'h3F;
		16'hC104: out_word = 8'hF1;
		16'hC105: out_word = 8'h18;
		16'hC106: out_word = 8'h0D;
		16'hC107: out_word = 8'h21;
		16'hC108: out_word = 8'hF8;
		16'hC109: out_word = 8'h5F;
		16'hC10A: out_word = 8'hF9;
		16'hC10B: out_word = 8'hEB;
		16'hC10C: out_word = 8'hD5;
		16'hC10D: out_word = 8'h21;
		16'hC10E: out_word = 8'h31;
		16'hC10F: out_word = 8'h3D;
		16'hC110: out_word = 8'h06;
		16'hC111: out_word = 8'h03;
		16'hC112: out_word = 8'hED;
		16'hC113: out_word = 8'hB0;
		16'hC114: out_word = 8'h08;
		16'hC115: out_word = 8'h21;
		16'hC116: out_word = 8'h47;
		16'hC117: out_word = 8'h01;
		16'hC118: out_word = 8'h11;
		16'hC119: out_word = 8'h07;
		16'hC11A: out_word = 8'h5C;
		16'hC11B: out_word = 8'h01;
		16'hC11C: out_word = 8'h1B;
		16'hC11D: out_word = 8'h00;
		16'hC11E: out_word = 8'hED;
		16'hC11F: out_word = 8'hB8;
		16'hC120: out_word = 8'hEB;
		16'hC121: out_word = 8'h23;
		16'hC122: out_word = 8'hDD;
		16'hC123: out_word = 8'h7D;
		16'hC124: out_word = 8'hFE;
		16'hC125: out_word = 8'h41;
		16'hC126: out_word = 8'h28;
		16'hC127: out_word = 8'h04;
		16'hC128: out_word = 8'h01;
		16'hC129: out_word = 8'h14;
		16'hC12A: out_word = 8'h00;
		16'hC12B: out_word = 8'h09;
		16'hC12C: out_word = 8'hE9;
		16'hC12D: out_word = 8'h01;
		16'hC12E: out_word = 8'hFD;
		16'hC12F: out_word = 8'h7F;
		16'hC130: out_word = 8'hAF;
		16'hC131: out_word = 8'hED;
		16'hC132: out_word = 8'h79;
		16'hC133: out_word = 8'h01;
		16'hC134: out_word = 8'hF7;
		16'hC135: out_word = 8'h3F;
		16'hC136: out_word = 8'h3E;
		16'hC137: out_word = 8'h81;
		16'hC138: out_word = 8'hED;
		16'hC139: out_word = 8'h79;
		16'hC13A: out_word = 8'h01;
		16'hC13B: out_word = 8'h77;
		16'hC13C: out_word = 8'hFF;
		16'hC13D: out_word = 8'h3E;
		16'hC13E: out_word = 8'hAB;
		16'hC13F: out_word = 8'hED;
		16'hC140: out_word = 8'h79;
		16'hC141: out_word = 8'h01;
		16'hC142: out_word = 8'hFD;
		16'hC143: out_word = 8'h7F;
		16'hC144: out_word = 8'h08;
		16'hC145: out_word = 8'hED;
		16'hC146: out_word = 8'h79;
		16'hC147: out_word = 8'hC9;
		16'hC148: out_word = 8'h01;
		16'hC149: out_word = 8'hFF;
		16'hC14A: out_word = 8'hFD;
		16'hC14B: out_word = 8'h7F;
		16'hC14C: out_word = 8'h3E;
		16'hC14D: out_word = 8'h10;
		16'hC14E: out_word = 8'hED;
		16'hC14F: out_word = 8'h79;
		16'hC150: out_word = 8'h21;
		16'hC151: out_word = 8'h0F;
		16'hC152: out_word = 8'hFF;
		16'hC153: out_word = 8'h01;
		16'hC154: out_word = 8'h22;
		16'hC155: out_word = 8'h09;
		16'hC156: out_word = 8'h5C;
		16'hC157: out_word = 8'hFB;
		16'hC158: out_word = 8'hCD;
		16'hC159: out_word = 8'h8E;
		16'hC15A: out_word = 8'h64;
		16'hC15B: out_word = 8'hFC;
		16'hC15C: out_word = 8'hDA;
		16'hC15D: out_word = 8'hC4;
		16'hC15E: out_word = 8'h61;
		16'hC15F: out_word = 8'h3E;
		16'hC160: out_word = 8'hFE;
		16'hC161: out_word = 8'hDB;
		16'hC162: out_word = 8'h6F;
		16'hC163: out_word = 8'hE6;
		16'hC164: out_word = 8'h08;
		16'hC165: out_word = 8'hCA;
		16'hC166: out_word = 8'h2C;
		16'hC167: out_word = 8'h34;
		16'hC168: out_word = 8'hF7;
		16'hC169: out_word = 8'hFD;
		16'hC16A: out_word = 8'hF7;
		16'hC16B: out_word = 8'hFE;
		16'hC16C: out_word = 8'h02;
		16'hC16D: out_word = 8'hC2;
		16'hC16E: out_word = 8'h16;
		16'hC16F: out_word = 8'h62;
		16'hC170: out_word = 8'h3A;
		16'hC171: out_word = 8'h95;
		16'hC172: out_word = 8'h60;
		16'hC173: out_word = 8'h04;
		16'hC174: out_word = 8'hFE;
		16'hC175: out_word = 8'h7F;
		16'hC176: out_word = 8'h26;
		16'hC177: out_word = 8'h21;
		16'hC178: out_word = 8'h27;
		16'hC179: out_word = 8'h65;
		16'hC17A: out_word = 8'hC3;
		16'hC17B: out_word = 8'h30;
		16'hC17C: out_word = 8'h0C;
		16'hC17D: out_word = 8'h87;
		16'hC17E: out_word = 8'hEB;
		16'hC17F: out_word = 8'h85;
		16'hC180: out_word = 8'h83;
		16'hC181: out_word = 8'h6F;
		16'hC182: out_word = 8'h01;
		16'hC183: out_word = 8'hF0;
		16'hC184: out_word = 8'h24;
		16'hC185: out_word = 8'h7E;
		16'hC186: out_word = 8'h23;
		16'hC187: out_word = 8'h66;
		16'hC188: out_word = 8'h7F;
		16'hC189: out_word = 8'hCD;
		16'hC18A: out_word = 8'h04;
		16'hC18B: out_word = 8'h62;
		16'hC18C: out_word = 8'h21;
		16'hC18D: out_word = 8'h0B;
		16'hC18E: out_word = 8'h65;
		16'hC18F: out_word = 8'h0A;
		16'hC190: out_word = 8'h07;
		16'hC191: out_word = 8'h17;
		16'hC192: out_word = 8'hFD;
		16'hC193: out_word = 8'hCB;
		16'hC194: out_word = 8'h01;
		16'hC195: out_word = 8'hFF;
		16'hC196: out_word = 8'hAE;
		16'hC197: out_word = 8'h76;
		16'hC198: out_word = 8'h21;
		16'hC199: out_word = 8'h03;
		16'hC19A: out_word = 8'h59;
		16'hC19B: out_word = 8'h36;
		16'hC19C: out_word = 8'h07;
		16'hC19D: out_word = 8'h2D;
		16'hC19E: out_word = 8'h72;
		16'hC19F: out_word = 8'hFD;
		16'hC1A0: out_word = 8'h05;
		16'hC1A1: out_word = 8'h9F;
		16'hC1A2: out_word = 8'hFD;
		16'hC1A3: out_word = 8'h11;
		16'hC1A4: out_word = 8'h04;
		16'hC1A5: out_word = 8'h59;
		16'hC1A6: out_word = 8'h01;
		16'hC1A7: out_word = 8'h7C;
		16'hC1A8: out_word = 8'hFF;
		16'hC1A9: out_word = 8'h00;
		16'hC1AA: out_word = 8'hED;
		16'hC1AB: out_word = 8'hB0;
		16'hC1AC: out_word = 8'h3E;
		16'hC1AD: out_word = 8'h38;
		16'hC1AE: out_word = 8'hCD;
		16'hC1AF: out_word = 8'hF8;
		16'hC1B0: out_word = 8'h60;
		16'hC1B1: out_word = 8'hF1;
		16'hC1B2: out_word = 8'h11;
		16'hC1B3: out_word = 8'h00;
		16'hC1B4: out_word = 8'h48;
		16'hC1B5: out_word = 8'h26;
		16'hC1B6: out_word = 8'h7C;
		16'hC1B7: out_word = 8'hE5;
		16'hC1B8: out_word = 8'hCD;
		16'hC1B9: out_word = 8'hAF;
		16'hC1BA: out_word = 8'h61;
		16'hC1BB: out_word = 8'h5F;
		16'hC1BC: out_word = 8'hFF;
		16'hC1BD: out_word = 8'h60;
		16'hC1BE: out_word = 8'hE1;
		16'hC1BF: out_word = 8'h24;
		16'hC1C0: out_word = 8'hFD;
		16'hC1C1: out_word = 8'hCB;
		16'hC1C2: out_word = 8'h74;
		16'hC1C3: out_word = 8'h28;
		16'hC1C4: out_word = 8'hF3;
		16'hC1C5: out_word = 8'h1E;
		16'hC1C6: out_word = 8'hA0;
		16'hC1C7: out_word = 8'hAA;
		16'hC1C8: out_word = 8'hEF;
		16'hC1C9: out_word = 8'h10;
		16'hC1CA: out_word = 8'h2B;
		16'hC1CB: out_word = 8'h42;
		16'hC1CC: out_word = 8'hEF;
		16'hC1CD: out_word = 8'h42;
		16'hC1CE: out_word = 8'hBD;
		16'hC1CF: out_word = 8'h6E;
		16'hC1D0: out_word = 8'hFF;
		16'hC1D1: out_word = 8'hBB;
		16'hC1D2: out_word = 8'h21;
		16'hC1D3: out_word = 8'h26;
		16'hC1D4: out_word = 8'h60;
		16'hC1D5: out_word = 8'hE5;
		16'hC1D6: out_word = 8'h2E;
		16'hC1D7: out_word = 8'h00;
		16'hC1D8: out_word = 8'h3A;
		16'hC1D9: out_word = 8'hF1;
		16'hC1DA: out_word = 8'h08;
		16'hC1DB: out_word = 8'h5C;
		16'hC1DC: out_word = 8'h2D;
		16'hC1DD: out_word = 8'hFE;
		16'hC1DE: out_word = 8'h38;
		16'hC1DF: out_word = 8'h28;
		16'hC1E0: out_word = 8'h41;
		16'hC1E1: out_word = 8'h2C;
		16'hC1E2: out_word = 8'h70;
		16'hC1E3: out_word = 8'h09;
		16'hC1E4: out_word = 8'hE2;
		16'hC1E5: out_word = 8'h3B;
		16'hC1E6: out_word = 8'h7C;
		16'hC1E7: out_word = 8'h0A;
		16'hC1E8: out_word = 8'h20;
		16'hC1E9: out_word = 8'h06;
		16'hC1EA: out_word = 8'h7D;
		16'hC1EB: out_word = 8'hC6;
		16'hC1EC: out_word = 8'h4F;
		16'hC1ED: out_word = 8'h6F;
		16'hC1EE: out_word = 8'h18;
		16'hC1EF: out_word = 8'h32;
		16'hC1F0: out_word = 8'hFE;
		16'hC1F1: out_word = 8'hA5;
		16'hC1F2: out_word = 8'h0B;
		16'hC1F3: out_word = 8'hF6;
		16'hC1F4: out_word = 8'hD6;
		16'hC1F5: out_word = 8'h3F;
		16'hC1F6: out_word = 8'hF6;
		16'hC1F7: out_word = 8'h28;
		16'hC1F8: out_word = 8'hCD;
		16'hC1F9: out_word = 8'hE6;
		16'hC1FA: out_word = 8'h60;
		16'hC1FB: out_word = 8'hD8;
		16'hC1FC: out_word = 8'h5F;
		16'hC1FD: out_word = 8'hE8;
		16'hC1FE: out_word = 8'h65;
		16'hC1FF: out_word = 8'hCB;
		16'hC200: out_word = 8'h3C;
		16'hC201: out_word = 8'hBF;
		16'hC202: out_word = 8'h1F;
		16'hC203: out_word = 8'h45;
		16'hC204: out_word = 8'h20;
		16'hC205: out_word = 8'h0C;
		16'hC206: out_word = 8'hC2;
		16'hC207: out_word = 8'hE6;
		16'hC208: out_word = 8'h0F;
		16'hC209: out_word = 8'hB4;
		16'hC20A: out_word = 8'h23;
		16'hC20B: out_word = 8'h7E;
		16'hC20C: out_word = 8'hFE;
		16'hC20D: out_word = 8'h18;
		16'hC20E: out_word = 8'h02;
		16'hC20F: out_word = 8'hE6;
		16'hC210: out_word = 8'hF0;
		16'hC211: out_word = 8'hB3;
		16'hC212: out_word = 8'hE5;
		16'hC213: out_word = 8'h92;
		16'hC214: out_word = 8'hE6;
		16'hC215: out_word = 8'h6F;
		16'hC216: out_word = 8'h34;
		16'hC217: out_word = 8'h60;
		16'hC218: out_word = 8'hA7;
		16'hC219: out_word = 8'h2C;
		16'hC21A: out_word = 8'h73;
		16'hC21B: out_word = 8'hBD;
		16'hC21C: out_word = 8'h7D;
		16'hC21D: out_word = 8'h32;
		16'hC21E: out_word = 8'h44;
		16'hC21F: out_word = 8'hC9;
		16'hC220: out_word = 8'hF9;
		16'hC221: out_word = 8'hF6;
		16'hC222: out_word = 8'h20;
		16'hC223: out_word = 8'hD6;
		16'hC224: out_word = 8'h30;
		16'hC225: out_word = 8'hD8;
		16'hC226: out_word = 8'hB8;
		16'hC227: out_word = 8'hC4;
		16'hC228: out_word = 8'h3F;
		16'hC229: out_word = 8'hD0;
		16'hC22A: out_word = 8'h83;
		16'hC22B: out_word = 8'h31;
		16'hC22C: out_word = 8'hD6;
		16'hC22D: out_word = 8'h87;
		16'hC22E: out_word = 8'h27;
		16'hC22F: out_word = 8'h10;
		16'hC230: out_word = 8'hE7;
		16'hC231: out_word = 8'h3F;
		16'hC232: out_word = 8'hC9;
		16'hC233: out_word = 8'h2A;
		16'hC234: out_word = 8'hEA;
		16'hC235: out_word = 8'h26;
		16'hC236: out_word = 8'h59;
		16'hC237: out_word = 8'h83;
		16'hC238: out_word = 8'h77;
		16'hC239: out_word = 8'hF5;
		16'hC23A: out_word = 8'hA7;
		16'hC23B: out_word = 8'h0F;
		16'hC23C: out_word = 8'hFF;
		16'hC23D: out_word = 8'hCD;
		16'hC23E: out_word = 8'h08;
		16'hC23F: out_word = 8'h61;
		16'hC240: out_word = 8'h94;
		16'hC241: out_word = 8'hF1;
		16'hC242: out_word = 8'hBE;
		16'hC243: out_word = 8'hE1;
		16'hC244: out_word = 8'hFF;
		16'hC245: out_word = 8'hCE;
		16'hC246: out_word = 8'h30;
		16'hC247: out_word = 8'h27;
		16'hC248: out_word = 8'hC5;
		16'hC249: out_word = 8'hD5;
		16'hC24A: out_word = 8'hE5;
		16'hC24B: out_word = 8'h87;
		16'hC24C: out_word = 8'hFE;
		16'hC24D: out_word = 8'h81;
		16'hC24E: out_word = 8'h40;
		16'hC24F: out_word = 8'h02;
		16'hC250: out_word = 8'hFC;
		16'hC251: out_word = 8'h3E;
		16'hC252: out_word = 8'h5C;
		16'hC253: out_word = 8'h6F;
		16'hC254: out_word = 8'h26;
		16'hC255: out_word = 8'h0F;
		16'hC256: out_word = 8'h29;
		16'hC257: out_word = 8'h7F;
		16'hC258: out_word = 8'h06;
		16'hC259: out_word = 8'h08;
		16'hC25A: out_word = 8'h7E;
		16'hC25B: out_word = 8'h12;
		16'hC25C: out_word = 8'hFF;
		16'hC25D: out_word = 8'h2C;
		16'hC25E: out_word = 8'h14;
		16'hC25F: out_word = 8'h10;
		16'hC260: out_word = 8'hFA;
		16'hC261: out_word = 8'hE1;
		16'hC262: out_word = 8'hD1;
		16'hC263: out_word = 8'hC1;
		16'hC264: out_word = 8'h1C;
		16'hC265: out_word = 8'hC8;
		16'hC266: out_word = 8'hC9;
		16'hC267: out_word = 8'hDD;
		16'hC268: out_word = 8'h67;
		16'hC269: out_word = 8'hBF;
		16'hC26A: out_word = 8'h7D;
		16'hC26B: out_word = 8'hD3;
		16'hC26C: out_word = 8'hFE;
		16'hC26D: out_word = 8'h11;
		16'hC26E: out_word = 8'h01;
		16'hC26F: out_word = 8'h8D;
		16'hC270: out_word = 8'h40;
		16'hC271: out_word = 8'h00;
		16'hC272: out_word = 8'hF9;
		16'hC273: out_word = 8'h06;
		16'hC274: out_word = 8'h62;
		16'hC275: out_word = 8'h69;
		16'hC276: out_word = 8'h36;
		16'hC277: out_word = 8'h7E;
		16'hC278: out_word = 8'h23;
		16'hC279: out_word = 8'h07;
		16'hC27A: out_word = 8'h02;
		16'hC27B: out_word = 8'h75;
		16'hC27C: out_word = 8'h4C;
		16'hC27D: out_word = 8'hFB;
		16'hC27E: out_word = 8'h08;
		16'hC27F: out_word = 8'h35;
		16'hC280: out_word = 8'hFF;
		16'hC281: out_word = 8'hFB;
		16'hC282: out_word = 8'h0E;
		16'hC283: out_word = 8'hAA;
		16'hC284: out_word = 8'h71;
		16'hC285: out_word = 8'h2C;
		16'hC286: out_word = 8'h20;
		16'hC287: out_word = 8'hFC;
		16'hC288: out_word = 8'h79;
		16'hC289: out_word = 8'hCF;
		16'hC28A: out_word = 8'h2F;
		16'hC28B: out_word = 8'h4F;
		16'hC28C: out_word = 8'h33;
		16'hC28D: out_word = 8'h5C;
		16'hC28E: out_word = 8'h28;
		16'hC28F: out_word = 8'hF4;
		16'hC290: out_word = 8'hF9;
		16'hC291: out_word = 8'h78;
		16'hC292: out_word = 8'hEE;
		16'hC293: out_word = 8'hC0;
		16'hC294: out_word = 8'h77;
		16'hC295: out_word = 8'h23;
		16'hC296: out_word = 8'hFE;
		16'hC297: out_word = 8'hE7;
		16'hC298: out_word = 8'h04;
		16'hC299: out_word = 8'hCB;
		16'hC29A: out_word = 8'h4C;
		16'hC29B: out_word = 8'hF4;
		16'hC29C: out_word = 8'h7D;
		16'hC29D: out_word = 8'hEE;
		16'hC29E: out_word = 8'hD0;
		16'hC29F: out_word = 8'h80;
		16'hC2A0: out_word = 8'h1F;
		16'hC2A1: out_word = 8'hF3;
		16'hC2A2: out_word = 8'hFF;
		16'hC2A3: out_word = 8'hE2;
		16'hC2A4: out_word = 8'hF6;
		16'hC2A5: out_word = 8'hFB;
		16'hC2A6: out_word = 8'h76;
		16'hC2A7: out_word = 8'hAF;
		16'hC2A8: out_word = 8'hDB;
		16'hC2A9: out_word = 8'hFE;
		16'hC2AA: out_word = 8'h2F;
		16'hC2AB: out_word = 8'hCF;
		16'hC2AC: out_word = 8'hE6;
		16'hC2AD: out_word = 8'h1F;
		16'hC2AE: out_word = 8'hF6;
		16'hC2AF: out_word = 8'hF3;
		16'hC2B0: out_word = 8'h9F;
		16'hC2B1: out_word = 8'h3C;
		16'hC2B2: out_word = 8'hE3;
		16'hC2B3: out_word = 8'hD3;
		16'hC2B4: out_word = 8'hFB;
		16'hC2B5: out_word = 8'h10;
		16'hC2B6: out_word = 8'h1F;
		16'hC2B7: out_word = 8'hFC;
		16'hC2B8: out_word = 8'h04;
		16'hC2B9: out_word = 8'h3D;
		16'hC2BA: out_word = 8'h20;
		16'hC2BB: out_word = 8'hFA;
		16'hC2BC: out_word = 8'h4F;
		16'hC2BD: out_word = 8'hEB;
		16'hC2BE: out_word = 8'h1F;
		16'hC2BF: out_word = 8'h38;
		16'hC2C0: out_word = 8'hEE;
		16'hC2C1: out_word = 8'hDD;
		16'hC2C2: out_word = 8'hFF;
		16'hC2C3: out_word = 8'h2C;
		16'hC2C4: out_word = 8'h18;
		16'hC2C5: out_word = 8'hA1;
		16'hC2C6: out_word = 8'hCD;
		16'hC2C7: out_word = 8'hA6;
		16'hC2C8: out_word = 8'h61;
		16'hC2C9: out_word = 8'h7C;
		16'hC2CA: out_word = 8'h01;
		16'hC2CB: out_word = 8'hF9;
		16'hC2CC: out_word = 8'hF7;
		16'hC2CD: out_word = 8'hDF;
		16'hC2CE: out_word = 8'hED;
		16'hC2CF: out_word = 8'h79;
		16'hC2D0: out_word = 8'h7D;
		16'hC2D1: out_word = 8'hFA;
		16'hC2D2: out_word = 8'h93;
		16'hC2D3: out_word = 8'hBF;
		16'hC2D4: out_word = 8'hFA;
		16'hC2D5: out_word = 8'hFB;
		16'hC2D6: out_word = 8'hEF;
		16'hC2D7: out_word = 8'hCF;
		16'hC2D8: out_word = 8'h3E;
		16'hC2D9: out_word = 8'h00;
		16'hC2DA: out_word = 8'hF9;
		16'hC2DB: out_word = 8'hFB;
		16'hC2DC: out_word = 8'hC9;
		16'hC2DD: out_word = 8'hF3;
		16'hC2DE: out_word = 8'h72;
		16'hC2DF: out_word = 8'hF6;
		16'hC2E0: out_word = 8'h80;
		16'hC2E1: out_word = 8'h6D;
		16'hC2E2: out_word = 8'hF6;
		16'hC2E3: out_word = 8'hC9;
		16'hC2E4: out_word = 8'hCE;
		16'hC2E5: out_word = 8'hDF;
		16'hC2E6: out_word = 8'h79;
		16'hC2E7: out_word = 8'hE0;
		16'hC2E8: out_word = 8'h78;
		16'hC2E9: out_word = 8'h67;
		16'hC2EA: out_word = 8'hCD;
		16'hC2EB: out_word = 8'h9D;
		16'hC2EC: out_word = 8'hF1;
		16'hC2ED: out_word = 8'hFA;
		16'hC2EE: out_word = 8'hA7;
		16'hC2EF: out_word = 8'hC9;
		16'hC2F0: out_word = 8'h21;
		16'hC2F1: out_word = 8'hA1;
		16'hC2F2: out_word = 8'h64;
		16'hC2F3: out_word = 8'hFF;
		16'hC2F4: out_word = 8'h77;
		16'hC2F5: out_word = 8'h76;
		16'hC2F6: out_word = 8'h01;
		16'hC2F7: out_word = 8'hFE;
		16'hC2F8: out_word = 8'h1F;
		16'hC2F9: out_word = 8'h21;
		16'hC2FA: out_word = 8'h60;
		16'hC2FB: out_word = 8'hFD;
		16'hC2FC: out_word = 8'h58;
		16'hC2FD: out_word = 8'hCD;
		16'hC2FE: out_word = 8'hDB;
		16'hC2FF: out_word = 8'h61;
		16'hC300: out_word = 8'h2E;
		16'hC301: out_word = 8'h09;
		16'hC302: out_word = 8'h3F;
		16'hC303: out_word = 8'hFB;
		16'hC304: out_word = 8'h18;
		16'hC305: out_word = 8'hEF;
		16'hC306: out_word = 8'h1E;
		16'hC307: out_word = 8'h04;
		16'hC308: out_word = 8'h16;
		16'hC309: out_word = 8'h05;
		16'hC30A: out_word = 8'h3F;
		16'hC30B: out_word = 8'hDC;
		16'hC30C: out_word = 8'h1F;
		16'hC30D: out_word = 8'h36;
		16'hC30E: out_word = 8'h07;
		16'hC30F: out_word = 8'h38;
		16'hC310: out_word = 8'h02;
		16'hC311: out_word = 8'h13;
		16'hC312: out_word = 8'h30;
		16'hC313: out_word = 8'h2C;
		16'hC314: out_word = 8'hFF;
		16'hC315: out_word = 8'h15;
		16'hC316: out_word = 8'h20;
		16'hC317: out_word = 8'hF5;
		16'hC318: out_word = 8'h7D;
		16'hC319: out_word = 8'hD6;
		16'hC31A: out_word = 8'h25;
		16'hC31B: out_word = 8'h6F;
		16'hC31C: out_word = 8'hCB;
		16'hC31D: out_word = 8'hF8;
		16'hC31E: out_word = 8'h00;
		16'hC31F: out_word = 8'h1D;
		16'hC320: out_word = 8'h20;
		16'hC321: out_word = 8'hE8;
		16'hC322: out_word = 8'h11;
		16'hC323: out_word = 8'hDF;
		16'hC324: out_word = 8'h61;
		16'hC325: out_word = 8'h1A;
		16'hC326: out_word = 8'hEE;
		16'hC327: out_word = 8'h01;
		16'hC328: out_word = 8'h12;
		16'hC329: out_word = 8'h06;
		16'hC32A: out_word = 8'hED;
		16'hC32B: out_word = 8'h90;
		16'hC32C: out_word = 8'hF9;
		16'hC32D: out_word = 8'h10;
		16'hC32E: out_word = 8'h60;
		16'hC32F: out_word = 8'hC9;
		16'hC330: out_word = 8'h7E;
		16'hC331: out_word = 8'h00;
		16'hC332: out_word = 8'h40;
		16'hC333: out_word = 8'h7E;
		16'hC334: out_word = 8'h23;
		16'hC335: out_word = 8'hB7;
		16'hC336: out_word = 8'hC8;
		16'hC337: out_word = 8'hBF;
		16'hC338: out_word = 8'h76;
		16'hC339: out_word = 8'h20;
		16'hC33A: out_word = 8'hFF;
		16'hC33B: out_word = 8'h04;
		16'hC33C: out_word = 8'h7A;
		16'hC33D: out_word = 8'hC6;
		16'hC33E: out_word = 8'h08;
		16'hC33F: out_word = 8'h57;
		16'hC340: out_word = 8'h18;
		16'hC341: out_word = 8'hF1;
		16'hC342: out_word = 8'h21;
		16'hC343: out_word = 8'hDD;
		16'hC344: out_word = 8'h11;
		16'hC345: out_word = 8'h66;
		16'hC346: out_word = 8'hFC;
		16'hC347: out_word = 8'h25;
		16'hC348: out_word = 8'h52;
		16'hC349: out_word = 8'h67;
		16'hC34A: out_word = 8'hF5;
		16'hC34B: out_word = 8'hE5;
		16'hC34C: out_word = 8'h5C;
		16'hC34D: out_word = 8'h01;
		16'hC34E: out_word = 8'h1E;
		16'hC34F: out_word = 8'hF1;
		16'hC350: out_word = 8'h3B;
		16'hC351: out_word = 8'h3A;
		16'hC352: out_word = 8'h36;
		16'hC353: out_word = 8'h0E;
		16'hC354: out_word = 8'h81;
		16'hC355: out_word = 8'h42;
		16'hC356: out_word = 8'hFA;
		16'hC357: out_word = 8'hC8;
		16'hC358: out_word = 8'hA4;
		16'hC359: out_word = 8'h07;
		16'hC35A: out_word = 8'hFA;
		16'hC35B: out_word = 8'hD6;
		16'hC35C: out_word = 8'h2A;
		16'hC35D: out_word = 8'h31;
		16'hC35E: out_word = 8'h42;
		16'hC35F: out_word = 8'hFA;
		16'hC360: out_word = 8'h0C;
		16'hC361: out_word = 8'hA4;
		16'hC362: out_word = 8'h14;
		16'hC363: out_word = 8'hFA;
		16'hC364: out_word = 8'h26;
		16'hC365: out_word = 8'h2A;
		16'hC366: out_word = 8'h25;
		16'hC367: out_word = 8'hFF;
		16'hC368: out_word = 8'h1D;
		16'hC369: out_word = 8'hC9;
		16'hC36A: out_word = 8'h32;
		16'hC36B: out_word = 8'hC2;
		16'hC36C: out_word = 8'hBB;
		16'hC36D: out_word = 8'h5C;
		16'hC36E: out_word = 8'hCF;
		16'hC36F: out_word = 8'hFD;
		16'hC370: out_word = 8'hFD;
		16'hC371: out_word = 8'h3C;
		16'hC372: out_word = 8'hFA;
		16'hC373: out_word = 8'h7F;
		16'hC374: out_word = 8'h42;
		16'hC375: out_word = 8'hD6;
		16'hC376: out_word = 8'h31;
		16'hC377: out_word = 8'hFF;
		16'hC378: out_word = 8'hFE;
		16'hC379: out_word = 8'h04;
		16'hC37A: out_word = 8'h30;
		16'hC37B: out_word = 8'hED;
		16'hC37C: out_word = 8'h0E;
		16'hC37D: out_word = 8'h01;
		16'hC37E: out_word = 8'hCD;
		16'hC37F: out_word = 8'h13;
		16'hC380: out_word = 8'h87;
		16'hC381: out_word = 8'h3D;
		16'hC382: out_word = 8'h18;
		16'hC383: out_word = 8'h49;
		16'hC384: out_word = 8'hFB;
		16'hC385: out_word = 8'hFD;
		16'hC386: out_word = 8'h7E;
		16'hC387: out_word = 8'hAF;
		16'hC388: out_word = 8'h00;
		16'hC389: out_word = 8'h7A;
		16'hC38A: out_word = 8'hA3;
		16'hC38B: out_word = 8'h21;
		16'hC38C: out_word = 8'hA4;
		16'hC38D: out_word = 8'h62;
		16'hC38E: out_word = 8'hE5;
		16'hC38F: out_word = 8'h7D;
		16'hC390: out_word = 8'h92;
		16'hC391: out_word = 8'hCD;
		16'hC392: out_word = 8'h68;
		16'hC393: out_word = 8'h64;
		16'hC394: out_word = 8'hD8;
		16'hC395: out_word = 8'h87;
		16'hC396: out_word = 8'h2E;
		16'hC397: out_word = 8'hFF;
		16'hC398: out_word = 8'h67;
		16'hC399: out_word = 8'h5E;
		16'hC39A: out_word = 8'hF7;
		16'hC39B: out_word = 8'h84;
		16'hC39C: out_word = 8'hFA;
		16'hC39D: out_word = 8'hFF;
		16'hC39E: out_word = 8'h6F;
		16'hC39F: out_word = 8'h22;
		16'hC3A0: out_word = 8'h92;
		16'hC3A1: out_word = 8'h62;
		16'hC3A2: out_word = 8'hEB;
		16'hC3A3: out_word = 8'hE1;
		16'hC3A4: out_word = 8'h01;
		16'hC3A5: out_word = 8'h05;
		16'hC3A6: out_word = 8'h1B;
		16'hC3A7: out_word = 8'h11;
		16'hC3A8: out_word = 8'hFF;
		16'hC3A9: out_word = 8'h1F;
		16'hC3AA: out_word = 8'h21;
		16'hC3AB: out_word = 8'h00;
		16'hC3AC: out_word = 8'hA2;
		16'hC3AD: out_word = 8'hA0;
		16'hC3AE: out_word = 8'hCD;
		16'hC3AF: out_word = 8'h1E;
		16'hC3B0: out_word = 8'hFA;
		16'hC3B1: out_word = 8'hD5;
		16'hC3B2: out_word = 8'hA2;
		16'hC3B3: out_word = 8'h06;
		16'hC3B4: out_word = 8'h01;
		16'hC3B5: out_word = 8'h7B;
		16'hC3B6: out_word = 8'hA1;
		16'hC3B7: out_word = 8'hCD;
		16'hC3B8: out_word = 8'h33;
		16'hC3B9: out_word = 8'h63;
		16'hC3BA: out_word = 8'h80;
		16'hC3BB: out_word = 8'hA3;
		16'hC3BC: out_word = 8'hF7;
		16'hC3BD: out_word = 8'h18;
		16'hC3BE: out_word = 8'h64;
		16'hC3BF: out_word = 8'h76;
		16'hC3C0: out_word = 8'hB9;
		16'hC3C1: out_word = 8'h9F;
		16'hC3C2: out_word = 8'hF6;
		16'hC3C3: out_word = 8'hCD;
		16'hC3C4: out_word = 8'h0C;
		16'hC3C5: out_word = 8'hB6;
		16'hC3C6: out_word = 8'h9E;
		16'hC3C7: out_word = 8'hA7;
		16'hC3C8: out_word = 8'hB6;
		16'hC3C9: out_word = 8'h2A;
		16'hC3CA: out_word = 8'h34;
		16'hC3CB: out_word = 8'h63;
		16'hC3CC: out_word = 8'h87;
		16'hC3CD: out_word = 8'h95;
		16'hC3CE: out_word = 8'h97;
		16'hC3CF: out_word = 8'h28;
		16'hC3D0: out_word = 8'h26;
		16'hC3D1: out_word = 8'h12;
		16'hC3D2: out_word = 8'h05;
		16'hC3D3: out_word = 8'h24;
		16'hC3D4: out_word = 8'h22;
		16'hC3D5: out_word = 8'h0F;
		16'hC3D6: out_word = 8'h08;
		16'hC3D7: out_word = 8'h20;
		16'hC3D8: out_word = 8'h03;
		16'hC3D9: out_word = 8'h2D;
		16'hC3DA: out_word = 8'hC1;
		16'hC3DB: out_word = 8'h18;
		16'hC3DC: out_word = 8'h1F;
		16'hC3DD: out_word = 8'h98;
		16'hC3DE: out_word = 8'h09;
		16'hC3DF: out_word = 8'hF9;
		16'hC3E0: out_word = 8'h2C;
		16'hC3E1: out_word = 8'h20;
		16'hC3E2: out_word = 8'h3F;
		16'hC3E3: out_word = 8'hC7;
		16'hC3E4: out_word = 8'hCB;
		16'hC3E5: out_word = 8'h34;
		16'hC3E6: out_word = 8'h6F;
		16'hC3E7: out_word = 8'h18;
		16'hC3E8: out_word = 8'hAF;
		16'hC3E9: out_word = 8'h0E;
		16'hC3EA: out_word = 8'h4A;
		16'hC3EB: out_word = 8'hCB;
		16'hC3EC: out_word = 8'h15;
		16'hC3ED: out_word = 8'h06;
		16'hC3EE: out_word = 8'h57;
		16'hC3EF: out_word = 8'hF6;
		16'hC3F0: out_word = 8'h04;
		16'hC3F1: out_word = 8'hC2;
		16'hC3F2: out_word = 8'h77;
		16'hC3F3: out_word = 8'h9E;
		16'hC3F4: out_word = 8'h3A;
		16'hC3F5: out_word = 8'hCC;
		16'hC3F6: out_word = 8'hAD;
		16'hC3F7: out_word = 8'h17;
		16'hC3F8: out_word = 8'h22;
		16'hC3F9: out_word = 8'h7F;
		16'hC3FA: out_word = 8'hFB;
		16'hC3FB: out_word = 8'hD0;
		16'hC3FC: out_word = 8'h18;
		16'hC3FD: out_word = 8'h38;
		16'hC3FE: out_word = 8'hFE;
		16'hC3FF: out_word = 8'h0C;
		16'hC400: out_word = 8'h20;
		16'hC401: out_word = 8'hE3;
		16'hC402: out_word = 8'h0E;
		16'hC403: out_word = 8'h2D;
		16'hC404: out_word = 8'h24;
		16'hC405: out_word = 8'hE3;
		16'hC406: out_word = 8'h7E;
		16'hC407: out_word = 8'h25;
		16'hC408: out_word = 8'hFF;
		16'hC409: out_word = 8'h77;
		16'hC40A: out_word = 8'hE5;
		16'hC40B: out_word = 8'hCD;
		16'hC40C: out_word = 8'hBA;
		16'hC40D: out_word = 8'h63;
		16'hC40E: out_word = 8'hE1;
		16'hC40F: out_word = 8'h18;
		16'hC410: out_word = 8'hFF;
		16'hC411: out_word = 8'hE3;
		16'hC412: out_word = 8'hFE;
		16'hC413: out_word = 8'hC7;
		16'hC414: out_word = 8'h20;
		16'hC415: out_word = 8'h10;
		16'hC416: out_word = 8'hE5;
		16'hC417: out_word = 8'h23;
		16'hC418: out_word = 8'h7E;
		16'hC419: out_word = 8'hC4;
		16'hC41A: out_word = 8'h2B;
		16'hC41B: out_word = 8'h77;
		16'hC41C: out_word = 8'hF9;
		16'hC41D: out_word = 8'h7C;
		16'hC41E: out_word = 8'hD6;
		16'hC41F: out_word = 8'hA1;
		16'hC420: out_word = 8'h20;
		16'hC421: out_word = 8'hF6;
		16'hC422: out_word = 8'hF8;
		16'hC423: out_word = 8'h3F;
		16'hC424: out_word = 8'hEC;
		16'hC425: out_word = 8'h12;
		16'hC426: out_word = 8'hFE;
		16'hC427: out_word = 8'hC9;
		16'hC428: out_word = 8'h20;
		16'hC429: out_word = 8'h1D;
		16'hC42A: out_word = 8'hCE;
		16'hC42B: out_word = 8'hE5;
		16'hC42C: out_word = 8'h4E;
		16'hC42D: out_word = 8'hEB;
		16'hC42E: out_word = 8'h71;
		16'hC42F: out_word = 8'h4F;
		16'hC430: out_word = 8'h69;
		16'hC431: out_word = 8'hEB;
		16'hC432: out_word = 8'h2B;
		16'hC433: out_word = 8'hEA;
		16'hC434: out_word = 8'hF5;
		16'hC435: out_word = 8'hA6;
		16'hC436: out_word = 8'hE1;
		16'hC437: out_word = 8'h67;
		16'hC438: out_word = 8'h7D;
		16'hC439: out_word = 8'hE6;
		16'hC43A: out_word = 8'h50;
		16'hC43B: out_word = 8'hB6;
		16'hC43C: out_word = 8'hCD;
		16'hC43D: out_word = 8'h1F;
		16'hC43E: out_word = 8'h87;
		16'hC43F: out_word = 8'h20;
		16'hC440: out_word = 8'hF9;
		16'hC441: out_word = 8'hC9;
		16'hC442: out_word = 8'hFC;
		16'hC443: out_word = 8'hFE;
		16'hC444: out_word = 8'h6C;
		16'hC445: out_word = 8'hD1;
		16'hC446: out_word = 8'hCA;
		16'hC447: out_word = 8'h6E;
		16'hC448: out_word = 8'h62;
		16'hC449: out_word = 8'h2F;
		16'hC44A: out_word = 8'h0D;
		16'hC44B: out_word = 8'h20;
		16'hC44C: out_word = 8'h09;
		16'hC44D: out_word = 8'hCD;
		16'hC44E: out_word = 8'hE7;
		16'hC44F: out_word = 8'h5A;
		16'hC450: out_word = 8'h1F;
		16'hC451: out_word = 8'h01;
		16'hC452: out_word = 8'h50;
		16'hC453: out_word = 8'hD2;
		16'hC454: out_word = 8'h91;
		16'hC455: out_word = 8'hFF;
		16'hC456: out_word = 8'h62;
		16'hC457: out_word = 8'hD5;
		16'hC458: out_word = 8'hCD;
		16'hC459: out_word = 8'hA8;
		16'hC45A: out_word = 8'h63;
		16'hC45B: out_word = 8'hD8;
		16'hC45C: out_word = 8'h4E;
		16'hC45D: out_word = 8'h17;
		16'hC45E: out_word = 8'h4E;
		16'hC45F: out_word = 8'hFF;
		16'hC460: out_word = 8'hAE;
		16'hC461: out_word = 8'hE6;
		16'hC462: out_word = 8'hF0;
		16'hC463: out_word = 8'h2E;
		16'hC464: out_word = 8'h77;
		16'hC465: out_word = 8'hC5;
		16'hC466: out_word = 8'hE7;
		16'hC467: out_word = 8'hA1;
		16'hC468: out_word = 8'hAF;
		16'hC469: out_word = 8'h32;
		16'hC46A: out_word = 8'h4C;
		16'hC46B: out_word = 8'hB3;
		16'hC46C: out_word = 8'h64;
		16'hC46D: out_word = 8'hDA;
		16'hC46E: out_word = 8'h3A;
		16'hC46F: out_word = 8'h3E;
		16'hC470: out_word = 8'hFF;
		16'hC471: out_word = 8'h01;
		16'hC472: out_word = 8'hEA;
		16'hC473: out_word = 8'h54;
		16'hC474: out_word = 8'hE8;
		16'hC475: out_word = 8'h1F;
		16'hC476: out_word = 8'h30;
		16'hC477: out_word = 8'h17;
		16'hC478: out_word = 8'h37;
		16'hC479: out_word = 8'h9E;
		16'hC47A: out_word = 8'hCB;
		16'hC47B: out_word = 8'h38;
		16'hC47C: out_word = 8'hD9;
		16'hC47D: out_word = 8'hE1;
		16'hC47E: out_word = 8'hC1;
		16'hC47F: out_word = 8'h62;
		16'hC480: out_word = 8'hCD;
		16'hC481: out_word = 8'h0F;
		16'hC482: out_word = 8'hB4;
		16'hC483: out_word = 8'h73;
		16'hC484: out_word = 8'h6F;
		16'hC485: out_word = 8'hC3;
		16'hC486: out_word = 8'hD5;
		16'hC487: out_word = 8'h62;
		16'hC488: out_word = 8'hF1;
		16'hC489: out_word = 8'h71;
		16'hC48A: out_word = 8'h79;
		16'hC48B: out_word = 8'hF5;
		16'hC48C: out_word = 8'h88;
		16'hC48D: out_word = 8'hF8;
		16'hC48E: out_word = 8'h3E;
		16'hC48F: out_word = 8'hE2;
		16'hC490: out_word = 8'h7C;
		16'hC491: out_word = 8'hF8;
		16'hC492: out_word = 8'h6F;
		16'hC493: out_word = 8'hD7;
		16'hC494: out_word = 8'h7F;
		16'hC495: out_word = 8'hBE;
		16'hC496: out_word = 8'h41;
		16'hC497: out_word = 8'h47;
		16'hC498: out_word = 8'h0E;
		16'hC499: out_word = 8'h03;
		16'hC49A: out_word = 8'hCD;
		16'hC49B: out_word = 8'hFD;
		16'hC49C: out_word = 8'h57;
		16'hC49D: out_word = 8'h74;
		16'hC49E: out_word = 8'h75;
		16'hC49F: out_word = 8'hA6;
		16'hC4A0: out_word = 8'h1C;
		16'hC4A1: out_word = 8'hE5;
		16'hC4A2: out_word = 8'hE4;
		16'hC4A3: out_word = 8'h50;
		16'hC4A4: out_word = 8'hF8;
		16'hC4A5: out_word = 8'h7B;
		16'hC4A6: out_word = 8'h2B;
		16'hC4A7: out_word = 8'hBE;
		16'hC4A8: out_word = 8'h28;
		16'hC4A9: out_word = 8'hC7;
		16'hC4AA: out_word = 8'h05;
		16'hC4AB: out_word = 8'h1D;
		16'hC4AC: out_word = 8'hFF;
		16'hC4AD: out_word = 8'hCD;
		16'hC4AE: out_word = 8'h53;
		16'hC4AF: out_word = 8'h64;
		16'hC4B0: out_word = 8'h23;
		16'hC4B1: out_word = 8'h10;
		16'hC4B2: out_word = 8'hEC;
		16'hC4B3: out_word = 8'hE1;
		16'hC4B4: out_word = 8'h1C;
		16'hC4B5: out_word = 8'h45;
		16'hC4B6: out_word = 8'hE8;
		16'hC4B7: out_word = 8'hF6;
		16'hC4B8: out_word = 8'h21;
		16'hC4B9: out_word = 8'hA9;
		16'hC4BA: out_word = 8'hE8;
		16'hC4BB: out_word = 8'h04;
		16'hC4BC: out_word = 8'hE9;
		16'hC4BD: out_word = 8'hA7;
		16'hC4BE: out_word = 8'h56;
		16'hC4BF: out_word = 8'hE9;
		16'hC4C0: out_word = 8'hED;
		16'hC4C1: out_word = 8'hC9;
		16'hC4C2: out_word = 8'hEB;
		16'hC4C3: out_word = 8'hAF;
		16'hC4C4: out_word = 8'h79;
		16'hC4C5: out_word = 8'hE9;
		16'hC4C6: out_word = 8'h7B;
		16'hC4C7: out_word = 8'h4F;
		16'hC4C8: out_word = 8'h78;
		16'hC4C9: out_word = 8'hFB;
		16'hC4CA: out_word = 8'hCD;
		16'hC4CB: out_word = 8'hFF;
		16'hC4CC: out_word = 8'hB0;
		16'hC4CD: out_word = 8'h22;
		16'hC4CE: out_word = 8'hEB;
		16'hC4CF: out_word = 8'hC9;
		16'hC4D0: out_word = 8'h3E;
		16'hC4D1: out_word = 8'h01;
		16'hC4D2: out_word = 8'h32;
		16'hC4D3: out_word = 8'h2A;
		16'hC4D4: out_word = 8'hC4;
		16'hC4D5: out_word = 8'h64;
		16'hC4D6: out_word = 8'h3A;
		16'hC4D7: out_word = 8'h17;
		16'hC4D8: out_word = 8'hB7;
		16'hC4D9: out_word = 8'hC8;
		16'hC4DA: out_word = 8'hDD;
		16'hC4DB: out_word = 8'h18;
		16'hC4DC: out_word = 8'h1B;
		16'hC4DD: out_word = 8'hF9;
		16'hC4DE: out_word = 8'hA3;
		16'hC4DF: out_word = 8'h7E;
		16'hC4E0: out_word = 8'hD0;
		16'hC4E1: out_word = 8'hFF;
		16'hC4E2: out_word = 8'hBE;
		16'hC4E3: out_word = 8'h3E;
		16'hC4E4: out_word = 8'h20;
		16'hC4E5: out_word = 8'h28;
		16'hC4E6: out_word = 8'h01;
		16'hC4E7: out_word = 8'h87;
		16'hC4E8: out_word = 8'h32;
		16'hC4E9: out_word = 8'h2C;
		16'hC4EA: out_word = 8'hCE;
		16'hC4EB: out_word = 8'h64;
		16'hC4EC: out_word = 8'hE1;
		16'hC4ED: out_word = 8'hE3;
		16'hC4EE: out_word = 8'hD6;
		16'hC4EF: out_word = 8'h20;
		16'hC4F0: out_word = 8'h90;
		16'hC4F1: out_word = 8'hE1;
		16'hC4F2: out_word = 8'hD0;
		16'hC4F3: out_word = 8'h30;
		16'hC4F4: out_word = 8'h00;
		16'hC4F5: out_word = 8'h2F;
		16'hC4F6: out_word = 8'h4A;
		16'hC4F7: out_word = 8'hDD;
		16'hC4F8: out_word = 8'hFE;
		16'hC4F9: out_word = 8'hB9;
		16'hC4FA: out_word = 8'h4F;
		16'hC4FB: out_word = 8'h1F;
		16'hC4FC: out_word = 8'h66;
		16'hC4FD: out_word = 8'hFF;
		16'hC4FE: out_word = 8'hE6;
		16'hC4FF: out_word = 8'h83;
		16'hC500: out_word = 8'h79;
		16'hC501: out_word = 8'h27;
		16'hC502: out_word = 8'h07;
		16'hC503: out_word = 8'h87;
		16'hC504: out_word = 8'hC6;
		16'hC505: out_word = 8'hD0;
		16'hC506: out_word = 8'h06;
		16'hC507: out_word = 8'h4F;
		16'hC508: out_word = 8'h7E;
		16'hC509: out_word = 8'hFC;
		16'hC50A: out_word = 8'h33;
		16'hC50B: out_word = 8'hB7;
		16'hC50C: out_word = 8'h20;
		16'hC50D: out_word = 8'h03;
		16'hC50E: out_word = 8'h1C;
		16'hC50F: out_word = 8'h18;
		16'hC510: out_word = 8'h54;
		16'hC511: out_word = 8'hA3;
		16'hC512: out_word = 8'hFF;
		16'hC513: out_word = 8'hC5;
		16'hC514: out_word = 8'hD5;
		16'hC515: out_word = 8'h06;
		16'hC516: out_word = 8'h04;
		16'hC517: out_word = 8'h1A;
		16'hC518: out_word = 8'h2F;
		16'hC519: out_word = 8'h12;
		16'hC51A: out_word = 8'h14;
		16'hC51B: out_word = 8'h73;
		16'hC51C: out_word = 8'hFC;
		16'hC51D: out_word = 8'h10;
		16'hC51E: out_word = 8'hF6;
		16'hC51F: out_word = 8'h77;
		16'hC520: out_word = 8'h4F;
		16'hC521: out_word = 8'hC4;
		16'hC522: out_word = 8'hEE;
		16'hC523: out_word = 8'h16;
		16'hC524: out_word = 8'h58;
		16'hC525: out_word = 8'h3E;
		16'hC526: out_word = 8'hD9;
		16'hC527: out_word = 8'hB0;
		16'hC528: out_word = 8'h12;
		16'hC529: out_word = 8'h1E;
		16'hC52A: out_word = 8'hDB;
		16'hC52B: out_word = 8'hE5;
		16'hC52C: out_word = 8'h3E;
		16'hC52D: out_word = 8'h07;
		16'hC52E: out_word = 8'h12;
		16'hC52F: out_word = 8'hE8;
		16'hC530: out_word = 8'hA3;
		16'hC531: out_word = 8'h0A;
		16'hC532: out_word = 8'hD8;
		16'hC533: out_word = 8'hF5;
		16'hC534: out_word = 8'h44;
		16'hC535: out_word = 8'hF8;
		16'hC536: out_word = 8'h61;
		16'hC537: out_word = 8'hDF;
		16'hC538: out_word = 8'hF1;
		16'hC539: out_word = 8'hC9;
		16'hC53A: out_word = 8'hDE;
		16'hC53B: out_word = 8'hA5;
		16'hC53C: out_word = 8'h18;
		16'hC53D: out_word = 8'h62;
		16'hC53E: out_word = 8'h69;
		16'hC53F: out_word = 8'hBB;
		16'hC540: out_word = 8'hAB;
		16'hC541: out_word = 8'h36;
		16'hC542: out_word = 8'hF3;
		16'hC543: out_word = 8'h07;
		16'hC544: out_word = 8'h01;
		16'hC545: out_word = 8'hFF;
		16'hC546: out_word = 8'h02;
		16'hC547: out_word = 8'hF9;
		16'hC548: out_word = 8'hC9;
		16'hC549: out_word = 8'hFF;
		16'hC54A: out_word = 8'h31;
		16'hC54B: out_word = 8'h32;
		16'hC54C: out_word = 8'h33;
		16'hC54D: out_word = 8'h34;
		16'hC54E: out_word = 8'h35;
		16'hC54F: out_word = 8'h36;
		16'hC550: out_word = 8'h37;
		16'hC551: out_word = 8'h38;
		16'hC552: out_word = 8'hEC;
		16'hC553: out_word = 8'h39;
		16'hC554: out_word = 8'h30;
		16'hC555: out_word = 8'h20;
		16'hC556: out_word = 8'h4D;
		16'hC557: out_word = 8'hFF;
		16'hC558: out_word = 8'h51;
		16'hC559: out_word = 8'hFF;
		16'hC55A: out_word = 8'h57;
		16'hC55B: out_word = 8'h45;
		16'hC55C: out_word = 8'h52;
		16'hC55D: out_word = 8'h54;
		16'hC55E: out_word = 8'h59;
		16'hC55F: out_word = 8'h55;
		16'hC560: out_word = 8'h49;
		16'hC561: out_word = 8'h4F;
		16'hC562: out_word = 8'hB1;
		16'hC563: out_word = 8'h50;
		16'hC564: out_word = 8'h47;
		16'hC565: out_word = 8'hE0;
		16'hC566: out_word = 8'h41;
		16'hC567: out_word = 8'h53;
		16'hC568: out_word = 8'h44;
		16'hC569: out_word = 8'hFE;
		16'hC56A: out_word = 8'h46;
		16'hC56B: out_word = 8'h47;
		16'hC56C: out_word = 8'h48;
		16'hC56D: out_word = 8'h4A;
		16'hC56E: out_word = 8'h4B;
		16'hC56F: out_word = 8'h4C;
		16'hC570: out_word = 8'h65;
		16'hC571: out_word = 8'hC5;
		16'hC572: out_word = 8'h1F;
		16'hC573: out_word = 8'hE0;
		16'hC574: out_word = 8'h63;
		16'hC575: out_word = 8'h5A;
		16'hC576: out_word = 8'h58;
		16'hC577: out_word = 8'h43;
		16'hC578: out_word = 8'h56;
		16'hC579: out_word = 8'hFD;
		16'hC57A: out_word = 8'h42;
		16'hC57B: out_word = 8'h4E;
		16'hC57C: out_word = 8'h4D;
		16'hC57D: out_word = 8'h73;
		16'hC57E: out_word = 8'h00;
		16'hC57F: out_word = 8'h20;
		16'hC580: out_word = 8'h8C;
		16'hC581: out_word = 8'hBD;
		16'hC582: out_word = 8'hFF;
		16'hC583: out_word = 8'h00;
		16'hC584: out_word = 8'h73;
		16'hC585: out_word = 8'h65;
		16'hC586: out_word = 8'h63;
		16'hC587: out_word = 8'hCE;
		16'hC588: out_word = 8'hFC;
		16'hC589: out_word = 8'h20;
		16'hC58A: out_word = 8'h61;
		16'hC58B: out_word = 8'h6C;
		16'hC58C: out_word = 8'h37;
		16'hC58D: out_word = 8'h72;
		16'hC58E: out_word = 8'h6D;
		16'hC58F: out_word = 8'h00;
		16'hC590: out_word = 8'h1B;
		16'hC591: out_word = 8'h69;
		16'hC592: out_word = 8'h6E;
		16'hC593: out_word = 8'h71;
		16'hC594: out_word = 8'hFC;
		16'hC595: out_word = 8'hAB;
		16'hC596: out_word = 8'hF2;
		16'hC597: out_word = 8'h68;
		16'hC598: out_word = 8'h6F;
		16'hC599: out_word = 8'h84;
		16'hC59A: out_word = 8'h75;
		16'hC59B: out_word = 8'hF3;
		16'hC59C: out_word = 8'hFB;
		16'hC59D: out_word = 8'h56;
		16'hC59E: out_word = 8'hF0;
		16'hC59F: out_word = 8'h5B;
		16'hC5A0: out_word = 8'h64;
		16'hC5A1: out_word = 8'h07;
		16'hC5A2: out_word = 8'h79;
		16'hC5A3: out_word = 8'h20;
		16'hC5A4: out_word = 8'h6F;
		16'hC5A5: out_word = 8'h8B;
		16'hC5A6: out_word = 8'h66;
		16'hC5A7: out_word = 8'h77;
		16'hC5A8: out_word = 8'h8F;
		16'hC5A9: out_word = 8'h65;
		16'hC5AA: out_word = 8'h6B;
		16'hC5AB: out_word = 8'hD0;
		16'hC5AC: out_word = 8'h5D;
		16'hC5AD: out_word = 8'h00;
		16'hC5AE: out_word = 8'hF3;
		16'hC5AF: out_word = 8'hF8;
		16'hC5B0: out_word = 8'hD4;
		16'hC5B1: out_word = 8'h6F;
		16'hC5B2: out_word = 8'h6E;
		16'hC5B3: out_word = 8'h74;
		16'hC5B4: out_word = 8'h68;
		16'hC5B5: out_word = 8'h40;
		16'hC5B6: out_word = 8'h48;
		16'hC5B7: out_word = 8'h65;
		16'hC5B8: out_word = 8'hE2;
		16'hC5B9: out_word = 8'h7C;
		16'hC5BA: out_word = 8'h23;
		16'hC5BB: out_word = 8'h32;
		16'hC5BC: out_word = 8'h30;
		16'hC5BD: out_word = 8'h48;
		16'hC5BE: out_word = 8'h62;
		16'hC5BF: out_word = 8'h9F;
		16'hC5C0: out_word = 8'h3D;
		16'hC5C1: out_word = 8'h6E;
		16'hC5C2: out_word = 8'h6F;
		16'hC5C3: out_word = 8'h42;
		16'hC5C4: out_word = 8'h43;
		16'hC5C5: out_word = 8'hFE;
		16'hC5C6: out_word = 8'h44;
		16'hC5C7: out_word = 8'h2C;
		16'hC5C8: out_word = 8'h62;
		16'hC5C9: out_word = 8'h31;
		16'hC5CA: out_word = 8'h3D;
		16'hC5CB: out_word = 8'h32;
		16'hC5CC: out_word = 8'h34;
		16'hC5CD: out_word = 8'hE1;
		16'hC5CE: out_word = 8'hC6;
		16'hC5CF: out_word = 8'hF6;
		16'hC5D0: out_word = 8'hE4;
		16'hC5D1: out_word = 8'h30;
		16'hC5D2: out_word = 8'h3D;
		16'hC5D3: out_word = 8'h73;
		16'hC5D4: out_word = 8'hE1;
		16'hC5D5: out_word = 8'h52;
		16'hC5D6: out_word = 8'hD8;
		16'hC5D7: out_word = 8'h67;
		16'hC5D8: out_word = 8'hC2;
		16'hC5D9: out_word = 8'h69;
		16'hC5DA: out_word = 8'hD4;
		16'hC5DB: out_word = 8'h20;
		16'hC5DC: out_word = 8'h62;
		16'hC5DD: out_word = 8'h0C;
		16'hC5DE: out_word = 8'h4C;
		16'hC5DF: out_word = 8'h73;
		16'hC5E0: out_word = 8'h5D;
		16'hC5E1: out_word = 8'h83;
		16'hC5E2: out_word = 8'hF5;
		16'hC5E3: out_word = 8'h37;
		16'hC5E4: out_word = 8'h8B;
		16'hC5E5: out_word = 8'h3D;
		16'hC5E6: out_word = 8'h61;
		16'hC5E7: out_word = 8'h8F;
		16'hC5E8: out_word = 8'h74;
		16'hC5E9: out_word = 8'h65;
		16'hC5EA: out_word = 8'h9F;
		16'hC5EB: out_word = 8'h72;
		16'hC5EC: out_word = 8'hB0;
		16'hC5ED: out_word = 8'h6C;
		16'hC5EE: out_word = 8'h6F;
		16'hC5EF: out_word = 8'h77;
		16'hC5F0: out_word = 8'h5D;
		16'hC5F1: out_word = 8'h31;
		16'hC5F2: out_word = 8'hB8;
		16'hC5F3: out_word = 8'h65;
		16'hC5F4: out_word = 8'hA6;
		16'hC5F5: out_word = 8'h20;
		16'hC5F6: out_word = 8'hB4;
		16'hC5F7: out_word = 8'h64;
		16'hC5F8: out_word = 8'h69;
		16'hC5F9: out_word = 8'h35;
		16'hC5FA: out_word = 8'h28;
		16'hC5FB: out_word = 8'hE6;
		16'hC5FC: out_word = 8'h73;
		16'hC5FD: out_word = 8'h49;
		16'hC5FE: out_word = 8'hED;
		16'hC5FF: out_word = 8'h29;
		16'hC600: out_word = 8'hA1;
		16'hC601: out_word = 8'hDE;
		16'hC602: out_word = 8'h72;
		16'hC603: out_word = 8'h76;
		16'hC604: out_word = 8'hF2;
		16'hC605: out_word = 8'h23;
		16'hC606: out_word = 8'h90;
		16'hC607: out_word = 8'hCC;
		16'hC608: out_word = 8'h29;
		16'hC609: out_word = 8'hA3;
		16'hC60A: out_word = 8'h41;
		16'hC60B: out_word = 8'h73;
		16'hC60C: out_word = 8'hFC;
		16'hC60D: out_word = 8'h34;
		16'hC60E: out_word = 8'h3E;
		16'hC60F: out_word = 8'hF3;
		16'hC610: out_word = 8'h6D;
		16'hC611: out_word = 8'h73;
		16'hC612: out_word = 8'h67;
		16'hC613: out_word = 8'h20;
		16'hC614: out_word = 8'h9D;
		16'hC615: out_word = 8'h61;
		16'hC616: out_word = 8'h66;
		16'hC617: out_word = 8'h6F;
		16'hC618: out_word = 8'h6C;
		16'hC619: out_word = 8'h09;
		16'hC61A: out_word = 8'hDC;
		16'hC61B: out_word = 8'hF7;
		16'hC61C: out_word = 8'hF3;
		16'hC61D: out_word = 8'h4C;
		16'hC61E: out_word = 8'hC7;
		16'hC61F: out_word = 8'h00;
		16'hC620: out_word = 8'h28;
		16'hC621: out_word = 8'h48;
		16'hC622: out_word = 8'h2C;
		16'hC623: out_word = 8'h50;
		16'hC624: out_word = 8'h36;
		16'hC625: out_word = 8'h21;
		16'hC626: out_word = 8'h3A;
		16'hC627: out_word = 8'h40;
		16'hC628: out_word = 8'h44;
		16'hC629: out_word = 8'h81;
		16'hC62A: out_word = 8'h49;
		16'hC62B: out_word = 8'h54;
		16'hC62C: out_word = 8'h02;
		16'hC62D: out_word = 8'h62;
		16'hC62E: out_word = 8'h04;
		16'hC62F: out_word = 8'h66;
		16'hC630: out_word = 8'h08;
		16'hC631: out_word = 8'h6C;
		16'hC632: out_word = 8'h10;
		16'hC633: out_word = 8'h71;
		16'hC634: out_word = 8'h20;
		16'hC635: out_word = 8'h75;
		16'hC636: out_word = 8'h40;
		16'hC637: out_word = 8'h92;
		16'hC638: out_word = 8'h81;
		16'hC639: out_word = 8'h9D;
		16'hC63A: out_word = 8'hAE;
		16'hC63B: out_word = 8'h02;
		16'hC63C: out_word = 8'h27;
		16'hC63D: out_word = 8'h04;
		16'hC63E: out_word = 8'hC1;
		16'hC63F: out_word = 8'h08;
		16'hC640: out_word = 8'hCE;
		16'hC641: out_word = 8'h10;
		16'hC642: out_word = 8'hD2;
		16'hC643: out_word = 8'h20;
		16'hC644: out_word = 8'h52;
		16'hC645: out_word = 8'h1E;
		16'hC646: out_word = 8'h78;
		16'hC647: out_word = 8'h74;
		16'hC648: out_word = 8'h2B;
		16'hC649: out_word = 8'h6B;
		16'hC64A: out_word = 8'h06;
		16'hC64B: out_word = 8'h79;
		16'hC64C: out_word = 8'h3A;
		16'hC64D: out_word = 8'hF7;
		16'hC64E: out_word = 8'h07;
		16'hC64F: out_word = 8'h53;
		16'hC650: out_word = 8'h70;
		16'hC651: out_word = 8'h61;
		16'hC652: out_word = 8'hFF;
		16'hC653: out_word = 8'h63;
		16'hC654: out_word = 8'h65;
		16'hC655: out_word = 8'h3D;
		16'hC656: out_word = 8'h54;
		16'hC657: out_word = 8'h52;
		16'hC658: out_word = 8'h44;
		16'hC659: out_word = 8'h4F;
		16'hC65A: out_word = 8'h53;
		16'hC65B: out_word = 8'h66;
		16'hC65C: out_word = 8'hFF;
		16'hC65D: out_word = 8'hED;
		16'hC65E: out_word = 8'h43;
		16'hC65F: out_word = 8'h53;
		16'hC660: out_word = 8'hCF;
		16'hC661: out_word = 8'h3D;
		16'hC662: out_word = 8'h42;
		16'hC663: out_word = 8'h4F;
		16'hC664: out_word = 8'h69;
		16'hC665: out_word = 8'h63;
		16'hC666: out_word = 8'h31;
		16'hC667: out_word = 8'hCB;
		16'hC668: out_word = 8'h32;
		16'hC669: out_word = 8'h38;
		16'hC66A: out_word = 8'hDA;
		16'hC66B: out_word = 8'h54;
		16'hC66C: out_word = 8'hF4;
		16'hC66D: out_word = 8'h34;
		16'hC66E: out_word = 8'hF9;
		16'hC66F: out_word = 8'hF5;
		16'hC670: out_word = 8'h44;
		16'hC671: out_word = 8'h3D;
		16'hC672: out_word = 8'h47;
		16'hC673: out_word = 8'h72;
		16'hC674: out_word = 8'hF5;
		16'hC675: out_word = 8'h1F;
		16'hC676: out_word = 8'h21;
		16'hC677: out_word = 8'h35;
		16'hC678: out_word = 8'h3F;
		16'hC679: out_word = 8'hE8;
		16'hC67A: out_word = 8'h62;
		16'hC67B: out_word = 8'h28;
		16'hC67C: out_word = 8'h50;
		16'hC67D: out_word = 8'h53;
		16'hC67E: out_word = 8'h42;
		16'hC67F: out_word = 8'hE8;
		16'hC680: out_word = 8'h5E;
		16'hC681: out_word = 8'h48;
		16'hC682: out_word = 8'h61;
		16'hC683: out_word = 8'h7B;
		16'hC684: out_word = 8'hBF;
		16'hC685: out_word = 8'hF5;
		16'hC686: out_word = 8'h6E;
		16'hC687: out_word = 8'h23;
		16'hC688: out_word = 8'hCE;
		16'hC689: out_word = 8'hF3;
		16'hC68A: out_word = 8'h30;
		16'hC68B: out_word = 8'h34;
		16'hC68C: out_word = 8'h29;
		16'hC68D: out_word = 8'hFA;
		16'hC68E: out_word = 8'h3D;
		16'hC68F: out_word = 8'h00;
		16'hC690: out_word = 8'h8D;
		16'hC691: out_word = 8'h69;
		16'hC692: out_word = 8'h72;
		16'hC693: out_word = 8'hE6;
		16'hC694: out_word = 8'h54;
		16'hC695: out_word = 8'h61;
		16'hC696: out_word = 8'h62;
		16'hC697: out_word = 8'h81;
		16'hC698: out_word = 8'h2B;
		16'hC699: out_word = 8'h21;
		16'hC69A: out_word = 8'hF7;
		16'hC69B: out_word = 8'h22;
		16'hC69C: out_word = 8'h32;
		16'hC69D: out_word = 8'hD3;
		16'hC69E: out_word = 8'h20;
		16'hC69F: out_word = 8'h91;
		16'hC6A0: out_word = 8'h73;
		16'hC6A1: out_word = 8'h2B;
		16'hC6A2: out_word = 8'hE3;
		16'hC6A3: out_word = 8'h43;
		16'hC6A4: out_word = 8'h4F;
		16'hC6A5: out_word = 8'h56;
		16'hC6A6: out_word = 8'h5B;
		16'hC6A7: out_word = 8'h58;
		16'hC6A8: out_word = 8'h89;
		16'hC6A9: out_word = 8'hA1;
		16'hC6AA: out_word = 8'hAC;
		16'hC6AB: out_word = 8'hD8;
		16'hC6AC: out_word = 8'hA0;
		16'hC6AD: out_word = 8'h4D;
		16'hC6AE: out_word = 8'h8B;
		16'hC6AF: out_word = 8'h27;
		16'hC6B0: out_word = 8'h72;
		16'hC6B1: out_word = 8'h55;
		16'hC6B2: out_word = 8'h70;
		16'hC6B3: out_word = 8'h09;
		16'hC6B4: out_word = 8'h85;
		16'hC6B5: out_word = 8'h29;
		16'hC6B6: out_word = 8'hFF;
		16'hC6B7: out_word = 8'h49;
		16'hC6B8: out_word = 8'h97;
		16'hC6B9: out_word = 8'hF3;
		16'hC6BA: out_word = 8'h47;
		16'hC6BB: out_word = 8'h6C;
		16'hC6BC: out_word = 8'h75;
		16'hC6BD: out_word = 8'h6B;
		16'hC6BE: out_word = 8'h0D;
		16'hC6BF: out_word = 8'h61;
		16'hC6C0: out_word = 8'h28;
		16'hC6C1: out_word = 8'h07;
		16'hC6C2: out_word = 8'h08;
		16'hC6C3: out_word = 8'h24;
		16'hC6C4: out_word = 8'h75;
		16'hC6C5: out_word = 8'hFF;
		16'hC6C6: out_word = 8'h37;
		16'hC6C7: out_word = 8'h31;
		16'hC6C8: out_word = 8'h2D;
		16'hC6C9: out_word = 8'h34;
		16'hC6CA: out_word = 8'h3D;
		16'hC6CB: out_word = 8'h64;
		16'hC6CC: out_word = 8'h72;
		16'hC6CD: out_word = 8'h69;
		16'hC6CE: out_word = 8'hE9;
		16'hC6CF: out_word = 8'h76;
		16'hC6D0: out_word = 8'h65;
		16'hC6D1: out_word = 8'h2C;
		16'hC6D2: out_word = 8'hE0;
		16'hC6D3: out_word = 8'h4D;
		16'hC6D4: out_word = 8'hAF;
		16'hC6D5: out_word = 8'h3D;
		16'hC6D6: out_word = 8'h9B;
		16'hC6D7: out_word = 8'hF3;
		16'hC6D8: out_word = 8'h89;
		16'hC6D9: out_word = 8'h79;
		16'hC6DA: out_word = 8'hFE;
		16'hC6DB: out_word = 8'hB7;
		16'hC6DC: out_word = 8'h70;
		16'hC6DD: out_word = 8'hEF;
		16'hC6DE: out_word = 8'h57;
		16'hC6DF: out_word = 8'h3D;
		16'hC6E0: out_word = 8'h75;
		16'hC6E1: out_word = 8'h6E;
		16'hC6E2: out_word = 8'h2F;
		16'hC6E3: out_word = 8'hFF;
		16'hC6E4: out_word = 8'hC3;
		16'hC6E5: out_word = 8'h20;
		16'hC6E6: out_word = 8'h74;
		16'hC6E7: out_word = 8'h75;
		16'hC6E8: out_word = 8'h72;
		16'hC6E9: out_word = 8'h29;
		16'hC6EA: out_word = 8'h72;
		16'hC6EB: out_word = 8'hE0;
		16'hC6EC: out_word = 8'h38;
		16'hC6ED: out_word = 8'h6C;
		16'hC6EE: out_word = 8'hEF;
		16'hC6EF: out_word = 8'h3A;
		16'hC6F0: out_word = 8'hE0;
		16'hC6F1: out_word = 8'h75;
		16'hC6F2: out_word = 8'h73;
		16'hC6F3: out_word = 8'h5B;
		16'hC6F4: out_word = 8'hDF;
		16'hC6F5: out_word = 8'h39;
		16'hC6F6: out_word = 8'hA5;
		16'hC6F7: out_word = 8'hDF;
		16'hC6F8: out_word = 8'h69;
		16'hC6F9: out_word = 8'hC7;
		16'hC6FA: out_word = 8'hA2;
		16'hC6FB: out_word = 8'h9D;
		16'hC6FC: out_word = 8'h26;
		16'hC6FD: out_word = 8'h0E;
		16'hC6FE: out_word = 8'h75;
		16'hC6FF: out_word = 8'h70;
		16'hC700: out_word = 8'h39;
		16'hC701: out_word = 8'h49;
		16'hC702: out_word = 8'h90;
		16'hC703: out_word = 8'h63;
		16'hC704: out_word = 8'h18;
		16'hC705: out_word = 8'hFC;
		16'hC706: out_word = 8'h64;
		16'hC707: out_word = 8'h20;
		16'hC708: out_word = 8'h6F;
		16'hC709: out_word = 8'h70;
		16'hC70A: out_word = 8'h97;
		16'hC70B: out_word = 8'hE7;
		16'hC70C: out_word = 8'hDE;
		16'hC70D: out_word = 8'hAE;
		16'hC70E: out_word = 8'h3D;
		16'hC70F: out_word = 8'h2E;
		16'hC710: out_word = 8'hF4;
		16'hC711: out_word = 8'hD6;
		16'hC712: out_word = 8'hFF;
		16'hC713: out_word = 8'h61;
		16'hC714: out_word = 8'h5E;
		16'hC715: out_word = 8'hFC;
		16'hC716: out_word = 8'h07;
		16'hC717: out_word = 8'h10;
		16'hC718: out_word = 8'h01;
		16'hC719: out_word = 8'h01;
		16'hC71A: out_word = 8'hC5;
		16'hC71B: out_word = 8'hFF;
		16'hC71C: out_word = 8'hA0;
		16'hC71D: out_word = 8'hD4;
		16'hC71E: out_word = 8'h25;
		16'hC71F: out_word = 8'h0B;
		16'hC720: out_word = 8'hFA;
		16'hC721: out_word = 8'hE9;
		16'hC722: out_word = 8'hF8;
		16'hC723: out_word = 8'h10;
		16'hC724: out_word = 8'hF1;
		16'hC725: out_word = 8'hCF;
		16'hC726: out_word = 8'h3C;
		16'hC727: out_word = 8'h40;
		16'hC728: out_word = 8'hE2;
		16'hC729: out_word = 8'hCC;
		16'hC72A: out_word = 8'h01;
		16'hC72B: out_word = 8'hFC;
		16'hC72C: out_word = 8'h84;
		16'hC72D: out_word = 8'h5F;
		16'hC72E: out_word = 8'hD9;
		16'hC72F: out_word = 8'hFF;
		16'hC730: out_word = 8'h07;
		16'hC731: out_word = 8'h39;
		16'hC732: out_word = 8'hFD;
		16'hC733: out_word = 8'h3B;
		16'hC734: out_word = 8'h5D;
		16'hC735: out_word = 8'hFC;
		16'hC736: out_word = 8'h88;
		16'hC737: out_word = 8'h26;
		16'hC738: out_word = 8'hE4;
		16'hC739: out_word = 8'hF8;
		16'hC73A: out_word = 8'h48;
		16'hC73B: out_word = 8'h28;
		16'hC73C: out_word = 8'h3A;
		16'hC73D: out_word = 8'h10;
		16'hC73E: out_word = 8'h3C;
		16'hC73F: out_word = 8'hA5;
		16'hC740: out_word = 8'h41;
		16'hC741: out_word = 8'hFC;
		16'hC742: out_word = 8'h20;
		16'hC743: out_word = 8'hF2;
		16'hC744: out_word = 8'h3E;
		16'hC745: out_word = 8'h50;
		16'hC746: out_word = 8'h4A;
		16'hC747: out_word = 8'hFE;
		16'hC748: out_word = 8'h0C;
		16'hC749: out_word = 8'h92;
		16'hC74A: out_word = 8'h5C;
		16'hC74B: out_word = 8'h58;
		16'hC74C: out_word = 8'h02;
		16'hC74D: out_word = 8'h6C;
		16'hC74E: out_word = 8'hC5;
		16'hC74F: out_word = 8'hFF;
		16'hC750: out_word = 8'h58;
		16'hC751: out_word = 8'h20;
		16'hC752: out_word = 8'hA0;
		16'hC753: out_word = 8'h21;
		16'hC754: out_word = 8'h5C;
		16'hC755: out_word = 8'h5B;
		16'hC756: out_word = 8'hF5;
		16'hC757: out_word = 8'hF1;
		16'hC758: out_word = 8'hE0;
		16'hC759: out_word = 8'h50;
		16'hC75A: out_word = 8'h21;
		16'hC75B: out_word = 8'h18;
		16'hC75C: out_word = 8'hBA;
		16'hC75D: out_word = 8'h17;
		16'hC75E: out_word = 8'h01;
		16'hC75F: out_word = 8'h07;
		16'hC760: out_word = 8'h31;
		16'hC761: out_word = 8'hB9;
		16'hC762: out_word = 8'hF6;
		16'hC763: out_word = 8'hFF;
		16'hC764: out_word = 8'hFF;
		16'hC765: out_word = 8'h5F;
		16'hC766: out_word = 8'h30;
		16'hC767: out_word = 8'hB0;
		16'hC768: out_word = 8'hF4;
		16'hC769: out_word = 8'hD1;
		16'hC76A: out_word = 8'hFF;
		16'hC76B: out_word = 8'h90;
		16'hC76C: out_word = 8'hED;
		16'hC76D: out_word = 8'h9B;
		16'hC76E: out_word = 8'h6E;
		16'hC76F: out_word = 8'h46;
		16'hC770: out_word = 8'h61;
		16'hC771: out_word = 8'h96;
		16'hC772: out_word = 8'h2A;
		16'hC773: out_word = 8'h43;
		16'hC774: out_word = 8'h24;
		16'hC775: out_word = 8'hD0;
		16'hC776: out_word = 8'hA3;
		16'hC777: out_word = 8'h08;
		16'hC778: out_word = 8'hFF;
		16'hC779: out_word = 8'h65;
		16'hC77A: out_word = 8'hF4;
		16'hC77B: out_word = 8'h09;
		16'hC77C: out_word = 8'hAA;
		16'hC77D: out_word = 8'hCB;
		16'hC77E: out_word = 8'hFD;
		16'hC77F: out_word = 8'h93;
		16'hC780: out_word = 8'h47;
		16'hC781: out_word = 8'hAA;
		16'hC782: out_word = 8'hFD;
		16'hC783: out_word = 8'hCB;
		16'hC784: out_word = 8'hD3;
		16'hC785: out_word = 8'h02;
		16'hC786: out_word = 8'hE7;
		16'hC787: out_word = 8'hF7;
		16'hC788: out_word = 8'hF4;
		16'hC789: out_word = 8'h09;
		16'hC78A: out_word = 8'hE7;
		16'hC78B: out_word = 8'hA8;
		16'hC78C: out_word = 8'h10;
		16'hC78D: out_word = 8'h4B;
		16'hC78E: out_word = 8'hFB;
		16'hC78F: out_word = 8'hC4;
		16'hC790: out_word = 8'h15;
		16'hC791: out_word = 8'hE6;
		16'hC792: out_word = 8'h53;
		16'hC793: out_word = 8'h81;
		16'hC794: out_word = 8'h0F;
		16'hC795: out_word = 8'hFB;
		16'hC796: out_word = 8'h52;
		16'hC797: out_word = 8'hE6;
		16'hC798: out_word = 8'hF6;
		16'hC799: out_word = 8'h50;
		16'hC79A: out_word = 8'h80;
		16'hC79B: out_word = 8'h3F;
		16'hC79C: out_word = 8'hEA;
		16'hC79D: out_word = 8'h3A;
		16'hC79E: out_word = 8'hF7;
		16'hC79F: out_word = 8'hB6;
		16'hC7A0: out_word = 8'h22;
		16'hC7A1: out_word = 8'h76;
		16'hC7A2: out_word = 8'hC9;
		16'hC7A3: out_word = 8'h22;
		16'hC7A4: out_word = 8'h0D;
		16'hC7A5: out_word = 8'h80;
		16'hC7A6: out_word = 8'h01;
		16'hC7A7: out_word = 8'hF3;
		16'hC7A8: out_word = 8'hFC;
		16'hC7A9: out_word = 8'hAF;
		16'hC7AA: out_word = 8'hCD;
		16'hC7AB: out_word = 8'h36;
		16'hC7AC: out_word = 8'h63;
		16'hC7AD: out_word = 8'h3E;
		16'hC7AE: out_word = 8'h10;
		16'hC7AF: out_word = 8'h31;
		16'hC7B0: out_word = 8'h43;
		16'hC7B1: out_word = 8'hFF;
		16'hC7B2: out_word = 8'hFD;
		16'hC7B3: out_word = 8'hCB;
		16'hC7B4: out_word = 8'h37;
		16'hC7B5: out_word = 8'h9E;
		16'hC7B6: out_word = 8'h21;
		16'hC7B7: out_word = 8'h60;
		16'hC7B8: out_word = 8'h6F;
		16'hC7B9: out_word = 8'h11;
		16'hC7BA: out_word = 8'hF1;
		16'hC7BB: out_word = 8'h00;
		16'hC7BC: out_word = 8'h5C;
		16'hC7BD: out_word = 8'h01;
		16'hC7BE: out_word = 8'h70;
		16'hC7BF: out_word = 8'hB8;
		16'hC7C0: out_word = 8'hED;
		16'hC7C1: out_word = 8'hB0;
		16'hC7C2: out_word = 8'h21;
		16'hC7C3: out_word = 8'h18;
		16'hC7C4: out_word = 8'h3E;
		16'hC7C5: out_word = 8'hE5;
		16'hC7C6: out_word = 8'h98;
		16'hC7C7: out_word = 8'h03;
		16'hC7C8: out_word = 8'h13;
		16'hC7C9: out_word = 8'h9E;
		16'hC7CA: out_word = 8'hED;
		16'hC7CB: out_word = 8'h73;
		16'hC7CC: out_word = 8'h3D;
		16'hC7CD: out_word = 8'h5C;
		16'hC7CE: out_word = 8'h7F;
		16'hC7CF: out_word = 8'hFC;
		16'hC7D0: out_word = 8'h64;
		16'hC7D1: out_word = 8'h60;
		16'hC7D2: out_word = 8'hCD;
		16'hC7D3: out_word = 8'h6F;
		16'hC7D4: out_word = 8'h7A;
		16'hC7D5: out_word = 8'hFB;
		16'hC7D6: out_word = 8'hF0;
		16'hC7D7: out_word = 8'h76;
		16'hC7D8: out_word = 8'hF3;
		16'hC7D9: out_word = 8'h26;
		16'hC7DA: out_word = 8'h00;
		16'hC7DB: out_word = 8'h06;
		16'hC7DC: out_word = 8'hFF;
		16'hC7DD: out_word = 8'h82;
		16'hC7DE: out_word = 8'h2C;
		16'hC7DF: out_word = 8'h21;
		16'hC7E0: out_word = 8'h55;
		16'hC7E1: out_word = 8'h6C;
		16'hC7E2: out_word = 8'h20;
		16'hC7E3: out_word = 8'h04;
		16'hC7E4: out_word = 8'hCB;
		16'hC7E5: out_word = 8'hE2;
		16'hC7E6: out_word = 8'h96;
		16'hC7E7: out_word = 8'h18;
		16'hC7E8: out_word = 8'h15;
		16'hC7E9: out_word = 8'h74;
		16'hC7EA: out_word = 8'hD6;
		16'hC7EB: out_word = 8'h26;
		16'hC7EC: out_word = 8'h11;
		16'hC7ED: out_word = 8'hEF;
		16'hC7EE: out_word = 8'hF1;
		16'hC7EF: out_word = 8'hFE;
		16'hC7F0: out_word = 8'h55;
		16'hC7F1: out_word = 8'h28;
		16'hC7F2: out_word = 8'h07;
		16'hC7F3: out_word = 8'h22;
		16'hC7F4: out_word = 8'hAA;
		16'hC7F5: out_word = 8'h78;
		16'hC7F6: out_word = 8'h03;
		16'hC7F7: out_word = 8'hCD;
		16'hC7F8: out_word = 8'h95;
		16'hC7F9: out_word = 8'h82;
		16'hC7FA: out_word = 8'hB8;
		16'hC7FB: out_word = 8'hAE;
		16'hC7FC: out_word = 8'h62;
		16'hC7FD: out_word = 8'h58;
		16'hC7FE: out_word = 8'hAA;
		16'hC7FF: out_word = 8'h63;
		16'hC800: out_word = 8'h53;
		16'hC801: out_word = 8'h46;
		16'hC802: out_word = 8'hFD;
		16'hC803: out_word = 8'hCE;
		16'hC804: out_word = 8'h0B;
		16'hC805: out_word = 8'h21;
		16'hC806: out_word = 8'hCC;
		16'hC807: out_word = 8'hFE;
		16'hC808: out_word = 8'h6F;
		16'hC809: out_word = 8'h22;
		16'hC80A: out_word = 8'h5F;
		16'hC80B: out_word = 8'h64;
		16'hC80C: out_word = 8'hF3;
		16'hC80D: out_word = 8'h31;
		16'hC80E: out_word = 8'h00;
		16'hC80F: out_word = 8'h3B;
		16'hC810: out_word = 8'h70;
		16'hC811: out_word = 8'h9B;
		16'hC812: out_word = 8'h13;
		16'hC813: out_word = 8'h03;
		16'hC814: out_word = 8'hFD;
		16'hC815: out_word = 8'hFB;
		16'hC816: out_word = 8'hF8;
		16'hC817: out_word = 8'h85;
		16'hC818: out_word = 8'hAF;
		16'hC819: out_word = 8'h32;
		16'hC81A: out_word = 8'h51;
		16'hC81B: out_word = 8'h6C;
		16'hC81C: out_word = 8'h3F;
		16'hC81D: out_word = 8'h7A;
		16'hC81E: out_word = 8'h62;
		16'hC81F: out_word = 8'hDD;
		16'hC820: out_word = 8'h21;
		16'hC821: out_word = 8'hA9;
		16'hC822: out_word = 8'h83;
		16'hC823: out_word = 8'h66;
		16'hC824: out_word = 8'hB2;
		16'hC825: out_word = 8'hE7;
		16'hC826: out_word = 8'h79;
		16'hC827: out_word = 8'hFB;
		16'hC828: out_word = 8'h3A;
		16'hC829: out_word = 8'hB1;
		16'hC82A: out_word = 8'hE6;
		16'hC82B: out_word = 8'h02;
		16'hC82C: out_word = 8'hFF;
		16'hC82D: out_word = 8'h28;
		16'hC82E: out_word = 8'h0A;
		16'hC82F: out_word = 8'h76;
		16'hC830: out_word = 8'h3E;
		16'hC831: out_word = 8'hFA;
		16'hC832: out_word = 8'hDB;
		16'hC833: out_word = 8'hDF;
		16'hC834: out_word = 8'h2F;
		16'hC835: out_word = 8'hFC;
		16'hC836: out_word = 8'hE6;
		16'hC837: out_word = 8'h07;
		16'hC838: out_word = 8'h20;
		16'hC839: out_word = 8'hF6;
		16'hC83A: out_word = 8'hCD;
		16'hC83B: out_word = 8'h7E;
		16'hC83C: out_word = 8'hE7;
		16'hC83D: out_word = 8'hDA;
		16'hC83E: out_word = 8'hEF;
		16'hC83F: out_word = 8'h7F;
		16'hC840: out_word = 8'h6F;
		16'hC841: out_word = 8'h01;
		16'hC842: out_word = 8'hAE;
		16'hC843: out_word = 8'hF8;
		16'hC844: out_word = 8'h18;
		16'hC845: out_word = 8'h37;
		16'hC846: out_word = 8'hCD;
		16'hC847: out_word = 8'h8C;
		16'hC848: out_word = 8'h80;
		16'hC849: out_word = 8'h7F;
		16'hC84A: out_word = 8'h2C;
		16'hC84B: out_word = 8'hDD;
		16'hC84C: out_word = 8'hCB;
		16'hC84D: out_word = 8'h08;
		16'hC84E: out_word = 8'h4E;
		16'hC84F: out_word = 8'hFF;
		16'hC850: out_word = 8'hF5;
		16'hC851: out_word = 8'hC4;
		16'hC852: out_word = 8'h5F;
		16'hC853: out_word = 8'h81;
		16'hC854: out_word = 8'hF1;
		16'hC855: out_word = 8'h20;
		16'hC856: out_word = 8'h21;
		16'hC857: out_word = 8'hDD;
		16'hC858: out_word = 8'hF3;
		16'hC859: out_word = 8'h7E;
		16'hC85A: out_word = 8'h10;
		16'hC85B: out_word = 8'h3D;
		16'hC85C: out_word = 8'h18;
		16'hC85D: out_word = 8'h8B;
		16'hC85E: out_word = 8'hFD;
		16'hC85F: out_word = 8'h36;
		16'hC860: out_word = 8'hEA;
		16'hC861: out_word = 8'h16;
		16'hC862: out_word = 8'h8A;
		16'hC863: out_word = 8'hEA;
		16'hC864: out_word = 8'h51;
		16'hC865: out_word = 8'h7C;
		16'hC866: out_word = 8'hEA;
		16'hC867: out_word = 8'h0B;
		16'hC868: out_word = 8'hAF;
		16'hC869: out_word = 8'hDD;
		16'hC86A: out_word = 8'h77;
		16'hC86B: out_word = 8'h0F;
		16'hC86C: out_word = 8'hC2;
		16'hC86D: out_word = 8'hFD;
		16'hC86E: out_word = 8'h12;
		16'hC86F: out_word = 8'hCE;
		16'hC870: out_word = 8'h36;
		16'hC871: out_word = 8'h13;
		16'hC872: out_word = 8'h5F;
		16'hC873: out_word = 8'hE2;
		16'hC874: out_word = 8'h7F;
		16'hC875: out_word = 8'h8E;
		16'hC876: out_word = 8'h81;
		16'hC877: out_word = 8'h3D;
		16'hC878: out_word = 8'hC3;
		16'hC879: out_word = 8'hA8;
		16'hC87A: out_word = 8'hCA;
		16'hC87B: out_word = 8'hE6;
		16'hC87C: out_word = 8'h3B;
		16'hC87D: out_word = 8'h61;
		16'hC87E: out_word = 8'h2A;
		16'hC87F: out_word = 8'h7B;
		16'hC880: out_word = 8'hE5;
		16'hC881: out_word = 8'h9F;
		16'hC882: out_word = 8'h71;
		16'hC883: out_word = 8'hC1;
		16'hC884: out_word = 8'hA7;
		16'hC885: out_word = 8'hED;
		16'hC886: out_word = 8'h42;
		16'hC887: out_word = 8'h28;
		16'hC888: out_word = 8'hF1;
		16'hC889: out_word = 8'h06;
		16'hC88A: out_word = 8'hCD;
		16'hC88B: out_word = 8'hF4;
		16'hC88C: out_word = 8'h86;
		16'hC88D: out_word = 8'h7F;
		16'hC88E: out_word = 8'h18;
		16'hC88F: out_word = 8'h64;
		16'hC890: out_word = 8'h01;
		16'hC891: out_word = 8'hDF;
		16'hC892: out_word = 8'hFA;
		16'hC893: out_word = 8'hED;
		16'hC894: out_word = 8'hCF;
		16'hC895: out_word = 8'h78;
		16'hC896: out_word = 8'hE6;
		16'hC897: out_word = 8'h4B;
		16'hC898: out_word = 8'h06;
		16'hC899: out_word = 8'h28;
		16'hC89A: out_word = 8'h12;
		16'hC89B: out_word = 8'h13;
		16'hC89C: out_word = 8'h05;
		16'hC89D: out_word = 8'hCA;
		16'hC89E: out_word = 8'h9C;
		16'hC89F: out_word = 8'h62;
		16'hC8A0: out_word = 8'h22;
		16'hC8A1: out_word = 8'hA7;
		16'hC8A2: out_word = 8'h82;
		16'hC8A3: out_word = 8'h87;
		16'hC8A4: out_word = 8'h22;
		16'hC8A5: out_word = 8'h94;
		16'hC8A6: out_word = 8'h39;
		16'hC8A7: out_word = 8'h89;
		16'hC8A8: out_word = 8'h5E;
		16'hC8A9: out_word = 8'h64;
		16'hC8AA: out_word = 8'h92;
		16'hC8AB: out_word = 8'h02;
		16'hC8AC: out_word = 8'hBF;
		16'hC8AD: out_word = 8'h1F;
		16'hC8AE: out_word = 8'hA7;
		16'hC8AF: out_word = 8'h28;
		16'hC8B0: out_word = 8'h08;
		16'hC8B1: out_word = 8'h8D;
		16'hC8B2: out_word = 8'h32;
		16'hC8B3: out_word = 8'h5C;
		16'hC8B4: out_word = 8'hFA;
		16'hC8B5: out_word = 8'hCD;
		16'hC8B6: out_word = 8'h71;
		16'hC8B7: out_word = 8'h63;
		16'hC8B8: out_word = 8'h18;
		16'hC8B9: out_word = 8'h2E;
		16'hC8BA: out_word = 8'h7F;
		16'hC8BB: out_word = 8'hD2;
		16'hC8BC: out_word = 8'h38;
		16'hC8BD: out_word = 8'h14;
		16'hC8BE: out_word = 8'h2A;
		16'hC8BF: out_word = 8'h6C;
		16'hC8C0: out_word = 8'h61;
		16'hC8C1: out_word = 8'h7C;
		16'hC8C2: out_word = 8'hB5;
		16'hC8C3: out_word = 8'hE3;
		16'hC8C4: out_word = 8'h28;
		16'hC8C5: out_word = 8'h5E;
		16'hC8C6: out_word = 8'hDD;
		16'hC8C7: out_word = 8'h7C;
		16'hC8C8: out_word = 8'h0F;
		16'hC8C9: out_word = 8'h16;
		16'hC8CA: out_word = 8'h00;
		16'hC8CB: out_word = 8'h19;
		16'hC8CC: out_word = 8'h11;
		16'hC8CD: out_word = 8'hFB;
		16'hC8CE: out_word = 8'hE6;
		16'hC8CF: out_word = 8'hED;
		16'hC8D0: out_word = 8'hA0;
		16'hC8D1: out_word = 8'h18;
		16'hC8D2: out_word = 8'h51;
		16'hC8D3: out_word = 8'hC9;
		16'hC8D4: out_word = 8'hCC;
		16'hC8D5: out_word = 8'h98;
		16'hC8D6: out_word = 8'h6E;
		16'hC8D7: out_word = 8'hF9;
		16'hC8D8: out_word = 8'hCC;
		16'hC8D9: out_word = 8'hAB;
		16'hC8DA: out_word = 8'h86;
		16'hC8DB: out_word = 8'hCA;
		16'hC8DC: out_word = 8'hD8;
		16'hC8DD: out_word = 8'hBD;
		16'hC8DE: out_word = 8'hE5;
		16'hC8DF: out_word = 8'h54;
		16'hC8E0: out_word = 8'h1F;
		16'hC8E1: out_word = 8'hD2;
		16'hC8E2: out_word = 8'hB7;
		16'hC8E3: out_word = 8'h27;
		16'hC8E4: out_word = 8'hA1;
		16'hC8E5: out_word = 8'h21;
		16'hC8E6: out_word = 8'hE1;
		16'hC8E7: out_word = 8'h7E;
		16'hC8E8: out_word = 8'h06;
		16'hC8E9: out_word = 8'h85;
		16'hC8EA: out_word = 8'h00;
		16'hC8EB: out_word = 8'h59;
		16'hC8EC: out_word = 8'hFF;
		16'hC8ED: out_word = 8'h6B;
		16'hC8EE: out_word = 8'h4E;
		16'hC8EF: out_word = 8'h51;
		16'hC8F0: out_word = 8'h23;
		16'hC8F1: out_word = 8'hED;
		16'hC8F2: out_word = 8'hB1;
		16'hC8F3: out_word = 8'h20;
		16'hC8F4: out_word = 8'h08;
		16'hC8F5: out_word = 8'hF9;
		16'hC8F6: out_word = 8'h21;
		16'hC8F7: out_word = 8'h65;
		16'hC8F8: out_word = 8'h6B;
		16'hC8F9: out_word = 8'h7A;
		16'hC8FA: out_word = 8'h91;
		16'hC8FB: out_word = 8'h4C;
		16'hC8FC: out_word = 8'h81;
		16'hC8FD: out_word = 8'h38;
		16'hC8FE: out_word = 8'h00;
		16'hC8FF: out_word = 8'h1E;
		16'hC900: out_word = 8'h4F;
		16'hC901: out_word = 8'h53;
		16'hC902: out_word = 8'hBB;
		16'hC903: out_word = 8'hD6;
		16'hC904: out_word = 8'h79;
		16'hC905: out_word = 8'hDD;
		16'hC906: out_word = 8'hF8;
		16'hC907: out_word = 8'h4E;
		16'hC908: out_word = 8'h02;
		16'hC909: out_word = 8'h5E;
		16'hC90A: out_word = 8'h23;
		16'hC90B: out_word = 8'h0D;
		16'hC90C: out_word = 8'hF2;
		16'hC90D: out_word = 8'h51;
		16'hC90E: out_word = 8'hDA;
		16'hC90F: out_word = 8'h94;
		16'hC910: out_word = 8'hE0;
		16'hC911: out_word = 8'h2B;
		16'hC912: out_word = 8'hE3;
		16'hC913: out_word = 8'h68;
		16'hC914: out_word = 8'h42;
		16'hC915: out_word = 8'h7A;
		16'hC916: out_word = 8'h50;
		16'hC917: out_word = 8'hC4;
		16'hC918: out_word = 8'h51;
		16'hC919: out_word = 8'h8C;
		16'hC91A: out_word = 8'h78;
		16'hC91B: out_word = 8'h09;
		16'hC91C: out_word = 8'h3E;
		16'hC91D: out_word = 8'h17;
		16'hC91E: out_word = 8'hEC;
		16'hC91F: out_word = 8'hC2;
		16'hC920: out_word = 8'h6E;
		16'hC921: out_word = 8'h06;
		16'hC922: out_word = 8'hFF;
		16'hC923: out_word = 8'h66;
		16'hC924: out_word = 8'h07;
		16'hC925: out_word = 8'h87;
		16'hC926: out_word = 8'h85;
		16'hC927: out_word = 8'h30;
		16'hC928: out_word = 8'h01;
		16'hC929: out_word = 8'h24;
		16'hC92A: out_word = 8'h6F;
		16'hC92B: out_word = 8'hE2;
		16'hC92C: out_word = 8'h7E;
		16'hC92D: out_word = 8'h23;
		16'hC92E: out_word = 8'h66;
		16'hC92F: out_word = 8'h7A;
		16'hC930: out_word = 8'hE9;
		16'hC931: out_word = 8'h08;
		16'hC932: out_word = 8'h7B;
		16'hC933: out_word = 8'h92;
		16'hC934: out_word = 8'h41;
		16'hC935: out_word = 8'hC0;
		16'hC936: out_word = 8'h4F;
		16'hC937: out_word = 8'h33;
		16'hC938: out_word = 8'hC9;
		16'hC939: out_word = 8'hC2;
		16'hC93A: out_word = 8'hF9;
		16'hC93B: out_word = 8'h7B;
		16'hC93C: out_word = 8'h4F;
		16'hC93D: out_word = 8'hAB;
		16'hC93E: out_word = 8'hDD;
		16'hC93F: out_word = 8'h21;
		16'hC940: out_word = 8'h53;
		16'hC941: out_word = 8'h6C;
		16'hC942: out_word = 8'hFD;
		16'hC943: out_word = 8'h35;
		16'hC944: out_word = 8'hF2;
		16'hC945: out_word = 8'hC9;
		16'hC946: out_word = 8'h61;
		16'hC947: out_word = 8'h36;
		16'hC948: out_word = 8'h02;
		16'hC949: out_word = 8'hCC;
		16'hC94A: out_word = 8'hC3;
		16'hC94B: out_word = 8'h04;
		16'hC94C: out_word = 8'hC8;
		16'hC94D: out_word = 8'h23;
		16'hC94E: out_word = 8'hF1;
		16'hC94F: out_word = 8'h6F;
		16'hC950: out_word = 8'h12;
		16'hC951: out_word = 8'h54;
		16'hC952: out_word = 8'h73;
		16'hC953: out_word = 8'hF6;
		16'hC954: out_word = 8'h10;
		16'hC955: out_word = 8'h07;
		16'hC956: out_word = 8'hFF;
		16'hC957: out_word = 8'hB5;
		16'hC958: out_word = 8'hFD;
		16'hC959: out_word = 8'h6F;
		16'hC95A: out_word = 8'h26;
		16'hC95B: out_word = 8'h0E;
		16'hC95C: out_word = 8'hCD;
		16'hC95D: out_word = 8'h13;
		16'hC95E: out_word = 8'h82;
		16'hC95F: out_word = 8'h1D;
		16'hC960: out_word = 8'hB2;
		16'hC961: out_word = 8'hF8;
		16'hC962: out_word = 8'h6B;
		16'hC963: out_word = 8'h6E;
		16'hC964: out_word = 8'hA8;
		16'hC965: out_word = 8'h24;
		16'hC966: out_word = 8'h92;
		16'hC967: out_word = 8'h2F;
		16'hC968: out_word = 8'hC3;
		16'hC969: out_word = 8'hC7;
		16'hC96A: out_word = 8'hF2;
		16'hC96B: out_word = 8'hD5;
		16'hC96C: out_word = 8'h3F;
		16'hC96D: out_word = 8'hB8;
		16'hC96E: out_word = 8'hFC;
		16'hC96F: out_word = 8'h44;
		16'hC970: out_word = 8'h2F;
		16'hC971: out_word = 8'h6F;
		16'hC972: out_word = 8'hF5;
		16'hC973: out_word = 8'hA7;
		16'hC974: out_word = 8'hF8;
		16'hC975: out_word = 8'hD9;
		16'hC976: out_word = 8'hF1;
		16'hC977: out_word = 8'hFE;
		16'hC978: out_word = 8'h55;
		16'hC979: out_word = 8'hFD;
		16'hC97A: out_word = 8'h21;
		16'hC97B: out_word = 8'h38;
		16'hC97C: out_word = 8'h6B;
		16'hC97D: out_word = 8'hCC;
		16'hC97E: out_word = 8'h5C;
		16'hC97F: out_word = 8'h7D;
		16'hC980: out_word = 8'h17;
		16'hC981: out_word = 8'hDF;
		16'hC982: out_word = 8'hFD;
		16'hC983: out_word = 8'h20;
		16'hC984: out_word = 8'h7E;
		16'hC985: out_word = 8'hEE;
		16'hC986: out_word = 8'h02;
		16'hC987: out_word = 8'h77;
		16'hC988: out_word = 8'h39;
		16'hC989: out_word = 8'h73;
		16'hC98A: out_word = 8'hAA;
		16'hC98B: out_word = 8'h63;
		16'hC98C: out_word = 8'hD4;
		16'hC98D: out_word = 8'hC1;
		16'hC98E: out_word = 8'h72;
		16'hC98F: out_word = 8'hEE;
		16'hC990: out_word = 8'h54;
		16'hC991: out_word = 8'h9E;
		16'hC992: out_word = 8'hEE;
		16'hC993: out_word = 8'h10;
		16'hC994: out_word = 8'h77;
		16'hC995: out_word = 8'h18;
		16'hC996: out_word = 8'h99;
		16'hC997: out_word = 8'hEF;
		16'hC998: out_word = 8'hBB;
		16'hC999: out_word = 8'hA8;
		16'hC99A: out_word = 8'hF7;
		16'hC99B: out_word = 8'hC3;
		16'hC99C: out_word = 8'h50;
		16'hC99D: out_word = 8'h1C;
		16'hC99E: out_word = 8'h02;
		16'hC99F: out_word = 8'h03;
		16'hC9A0: out_word = 8'hDA;
		16'hC9A1: out_word = 8'h20;
		16'hC9A2: out_word = 8'h15;
		16'hC9A3: out_word = 8'h7E;
		16'hC9A4: out_word = 8'h41;
		16'hC9A5: out_word = 8'hEF;
		16'hC9A6: out_word = 8'hEF;
		16'hC9A7: out_word = 8'hC1;
		16'hC9A8: out_word = 8'h42;
		16'hC9A9: out_word = 8'hBA;
		16'hC9AA: out_word = 8'hD0;
		16'hC9AB: out_word = 8'hE8;
		16'hC9AC: out_word = 8'h08;
		16'hC9AD: out_word = 8'h9C;
		16'hC9AE: out_word = 8'h4F;
		16'hC9AF: out_word = 8'h1F;
		16'hC9B0: out_word = 8'hC9;
		16'hC9B1: out_word = 8'hFD;
		16'hC9B2: out_word = 8'h7E;
		16'hC9B3: out_word = 8'hF8;
		16'hC9B4: out_word = 8'hCE;
		16'hC9B5: out_word = 8'hFE;
		16'hC9B6: out_word = 8'h0D;
		16'hC9B7: out_word = 8'hC8;
		16'hC9B8: out_word = 8'h37;
		16'hC9B9: out_word = 8'h1F;
		16'hC9BA: out_word = 8'h3A;
		16'hC9BB: out_word = 8'hF8;
		16'hC9BC: out_word = 8'h5C;
		16'hC9BD: out_word = 8'hC6;
		16'hC9BE: out_word = 8'h41;
		16'hC9BF: out_word = 8'hF8;
		16'hC9C0: out_word = 8'h32;
		16'hC9C1: out_word = 8'hE9;
		16'hC9C2: out_word = 8'h6A;
		16'hC9C3: out_word = 8'h21;
		16'hC9C4: out_word = 8'hD3;
		16'hC9C5: out_word = 8'hB2;
		16'hC9C6: out_word = 8'hC3;
		16'hC9C7: out_word = 8'hA4;
		16'hC9C8: out_word = 8'h14;
		16'hC9C9: out_word = 8'hEB;
		16'hC9CA: out_word = 8'h2A;
		16'hC9CB: out_word = 8'hCD;
		16'hC9CC: out_word = 8'h69;
		16'hC9CD: out_word = 8'hFA;
		16'hC9CE: out_word = 8'h04;
		16'hC9CF: out_word = 8'h6B;
		16'hC9D0: out_word = 8'hF4;
		16'hC9D1: out_word = 8'h3E;
		16'hC9D2: out_word = 8'hFE;
		16'hC9D3: out_word = 8'h07;
		16'hC9D4: out_word = 8'hCD;
		16'hC9D5: out_word = 8'hA1;
		16'hC9D6: out_word = 8'h7A;
		16'hC9D7: out_word = 8'h21;
		16'hC9D8: out_word = 8'hAC;
		16'hC9D9: out_word = 8'h69;
		16'hC9DA: out_word = 8'h82;
		16'hC9DB: out_word = 8'hEF;
		16'hC9DC: out_word = 8'hDC;
		16'hC9DD: out_word = 8'h60;
		16'hC9DE: out_word = 8'h60;
		16'hC9DF: out_word = 8'hF4;
		16'hC9E0: out_word = 8'hAF;
		16'hC9E1: out_word = 8'hC3;
		16'hC9E2: out_word = 8'h61;
		16'hC9E3: out_word = 8'h86;
		16'hC9E4: out_word = 8'h40;
		16'hC9E5: out_word = 8'hFE;
		16'hC9E6: out_word = 8'hA7;
		16'hC9E7: out_word = 8'hCA;
		16'hC9E8: out_word = 8'h33;
		16'hC9E9: out_word = 8'h63;
		16'hC9EA: out_word = 8'h3D;
		16'hC9EB: out_word = 8'h28;
		16'hC9EC: out_word = 8'h0D;
		16'hC9ED: out_word = 8'hF6;
		16'hC9EE: out_word = 8'h3A;
		16'hC9EF: out_word = 8'hC6;
		16'hC9F0: out_word = 8'h04;
		16'hC9F1: out_word = 8'hBD;
		16'hC9F2: out_word = 8'hC7;
		16'hC9F3: out_word = 8'hC3;
		16'hC9F4: out_word = 8'h9F;
		16'hC9F5: out_word = 8'h3C;
		16'hC9F6: out_word = 8'h3F;
		16'hC9F7: out_word = 8'h99;
		16'hC9F8: out_word = 8'h62;
		16'hC9F9: out_word = 8'h3E;
		16'hC9FA: out_word = 8'h30;
		16'hC9FB: out_word = 8'h00;
		16'hC9FC: out_word = 8'h50;
		16'hC9FD: out_word = 8'h0A;
		16'hC9FE: out_word = 8'h2F;
		16'hC9FF: out_word = 8'h73;
		16'hCA00: out_word = 8'h4E;
		16'hCA01: out_word = 8'hE6;
		16'hCA02: out_word = 8'h80;
		16'hCA03: out_word = 8'h0F;
		16'hCA04: out_word = 8'hFF;
		16'hCA05: out_word = 8'h32;
		16'hCA06: out_word = 8'h3C;
		16'hCA07: out_word = 8'hE1;
		16'hCA08: out_word = 8'h7D;
		16'hCA09: out_word = 8'hE6;
		16'hCA0A: out_word = 8'h03;
		16'hCA0B: out_word = 8'h22;
		16'hCA0C: out_word = 8'hD1;
		16'hCA0D: out_word = 8'hF7;
		16'hCA0E: out_word = 8'hD8;
		16'hCA0F: out_word = 8'h11;
		16'hCA10: out_word = 8'h20;
		16'hCA11: out_word = 8'h6E;
		16'hCA12: out_word = 8'hC3;
		16'hCA13: out_word = 8'h28;
		16'hCA14: out_word = 8'h03;
		16'hCA15: out_word = 8'h8F;
		16'hCA16: out_word = 8'h66;
		16'hCA17: out_word = 8'h21;
		16'hCA18: out_word = 8'hFB;
		16'hCA19: out_word = 8'h01;
		16'hCA1A: out_word = 8'h6B;
		16'hCA1B: out_word = 8'h72;
		16'hCA1C: out_word = 8'h23;
		16'hCA1D: out_word = 8'h73;
		16'hCA1E: out_word = 8'h98;
		16'hCA1F: out_word = 8'hBB;
		16'hCA20: out_word = 8'h21;
		16'hCA21: out_word = 8'h47;
		16'hCA22: out_word = 8'h98;
		16'hCA23: out_word = 8'h28;
		16'hCA24: out_word = 8'h09;
		16'hCA25: out_word = 8'h70;
		16'hCA26: out_word = 8'h4D;
		16'hCA27: out_word = 8'hE4;
		16'hCA28: out_word = 8'h3D;
		16'hCA29: out_word = 8'hE8;
		16'hCA2A: out_word = 8'h28;
		16'hCA2B: out_word = 8'h4A;
		16'hCA2C: out_word = 8'h5E;
		16'hCA2D: out_word = 8'h11;
		16'hCA2E: out_word = 8'h19;
		16'hCA2F: out_word = 8'h6B;
		16'hCA30: out_word = 8'h0E;
		16'hCA31: out_word = 8'h06;
		16'hCA32: out_word = 8'hED;
		16'hCA33: out_word = 8'hB0;
		16'hCA34: out_word = 8'hD3;
		16'hCA35: out_word = 8'hFF;
		16'hCA36: out_word = 8'hDC;
		16'hCA37: out_word = 8'h11;
		16'hCA38: out_word = 8'h09;
		16'hCA39: out_word = 8'h6A;
		16'hCA3A: out_word = 8'h2E;
		16'hCA3B: out_word = 8'h00;
		16'hCA3C: out_word = 8'h8B;
		16'hCA3D: out_word = 8'hCD;
		16'hCA3E: out_word = 8'h82;
		16'hCA3F: out_word = 8'h02;
		16'hCA40: out_word = 8'h3A;
		16'hCA41: out_word = 8'h72;
		16'hCA42: out_word = 8'hF8;
		16'hCA43: out_word = 8'h01;
		16'hCA44: out_word = 8'hC3;
		16'hCA45: out_word = 8'hF8;
		16'hCA46: out_word = 8'hDF;
		16'hCA47: out_word = 8'hCD;
		16'hCA48: out_word = 8'h0B;
		16'hCA49: out_word = 8'h5E;
		16'hCA4A: out_word = 8'hDF;
		16'hCA4B: out_word = 8'h28;
		16'hCA4C: out_word = 8'h0A;
		16'hCA4D: out_word = 8'h26;
		16'hCA4E: out_word = 8'h10;
		16'hCA4F: out_word = 8'h89;
		16'hCA50: out_word = 8'h99;
		16'hCA51: out_word = 8'hA2;
		16'hCA52: out_word = 8'h50;
		16'hCA53: out_word = 8'h24;
		16'hCA54: out_word = 8'hA2;
		16'hCA55: out_word = 8'hFD;
		16'hCA56: out_word = 8'h2C;
		16'hCA57: out_word = 8'h19;
		16'hCA58: out_word = 8'h5D;
		16'hCA59: out_word = 8'h5F;
		16'hCA5A: out_word = 8'hF6;
		16'hCA5B: out_word = 8'h5C;
		16'hCA5C: out_word = 8'h6F;
		16'hCA5D: out_word = 8'h67;
		16'hCA5E: out_word = 8'h90;
		16'hCA5F: out_word = 8'h22;
		16'hCA60: out_word = 8'h36;
		16'hCA61: out_word = 8'h7E;
		16'hCA62: out_word = 8'h3C;
		16'hCA63: out_word = 8'h32;
		16'hCA64: out_word = 8'h16;
		16'hCA65: out_word = 8'h5D;
		16'hCA66: out_word = 8'hC9;
		16'hCA67: out_word = 8'h9F;
		16'hCA68: out_word = 8'h8E;
		16'hCA69: out_word = 8'h01;
		16'hCA6A: out_word = 8'hF7;
		16'hCA6B: out_word = 8'hEF;
		16'hCA6C: out_word = 8'hED;
		16'hCA6D: out_word = 8'h79;
		16'hCA6E: out_word = 8'hFE;
		16'hCA6F: out_word = 8'hC9;
		16'hCA70: out_word = 8'h3E;
		16'hCA71: out_word = 8'h10;
		16'hCA72: out_word = 8'hC5;
		16'hCA73: out_word = 8'h01;
		16'hCA74: out_word = 8'hFD;
		16'hCA75: out_word = 8'h7F;
		16'hCA76: out_word = 8'h7F;
		16'hCA77: out_word = 8'hF7;
		16'hCA78: out_word = 8'hC1;
		16'hCA79: out_word = 8'hC9;
		16'hCA7A: out_word = 8'h21;
		16'hCA7B: out_word = 8'h8B;
		16'hCA7C: out_word = 8'h6C;
		16'hCA7D: out_word = 8'h3E;
		16'hCA7E: out_word = 8'h99;
		16'hCA7F: out_word = 8'h0D;
		16'hCA80: out_word = 8'hF4;
		16'hCA81: out_word = 8'hFF;
		16'hCA82: out_word = 8'hF4;
		16'hCA83: out_word = 8'hC4;
		16'hCA84: out_word = 8'h06;
		16'hCA85: out_word = 8'hBF;
		16'hCA86: out_word = 8'hFC;
		16'hCA87: out_word = 8'hAB;
		16'hCA88: out_word = 8'hD6;
		16'hCA89: out_word = 8'h01;
		16'hCA8A: out_word = 8'h30;
		16'hCA8B: out_word = 8'hF3;
		16'hCA8C: out_word = 8'hC9;
		16'hCA8D: out_word = 8'hFF;
		16'hCA8E: out_word = 8'hAD;
		16'hCA8F: out_word = 8'h0E;
		16'hCA90: out_word = 8'h15;
		16'hCA91: out_word = 8'h62;
		16'hCA92: out_word = 8'h6B;
		16'hCA93: out_word = 8'hCD;
		16'hCA94: out_word = 8'h67;
		16'hCA95: out_word = 8'h63;
		16'hCA96: out_word = 8'hFB;
		16'hCA97: out_word = 8'h20;
		16'hCA98: out_word = 8'hF8;
		16'hCA99: out_word = 8'h21;
		16'hCA9A: out_word = 8'h3F;
		16'hCA9B: out_word = 8'h07;
		16'hCA9C: out_word = 8'h94;
		16'hCA9D: out_word = 8'hE4;
		16'hCA9E: out_word = 8'h61;
		16'hCA9F: out_word = 8'hE4;
		16'hCAA0: out_word = 8'hD7;
		16'hCAA1: out_word = 8'h69;
		16'hCAA2: out_word = 8'hC9;
		16'hCAA3: out_word = 8'hDB;
		16'hCAA4: out_word = 8'hC8;
		16'hCAA5: out_word = 8'h7B;
		16'hCAA6: out_word = 8'h18;
		16'hCAA7: out_word = 8'hF4;
		16'hCAA8: out_word = 8'hC9;
		16'hCAA9: out_word = 8'hFF;
		16'hCAAA: out_word = 8'h2A;
		16'hCAAB: out_word = 8'h95;
		16'hCAAC: out_word = 8'h63;
		16'hCAAD: out_word = 8'h11;
		16'hCAAE: out_word = 8'h80;
		16'hCAAF: out_word = 8'hF7;
		16'hCAB0: out_word = 8'h06;
		16'hCAB1: out_word = 8'h08;
		16'hCAB2: out_word = 8'hF4;
		16'hCAB3: out_word = 8'h7E;
		16'hCAB4: out_word = 8'h12;
		16'hCAB5: out_word = 8'h13;
		16'hCAB6: out_word = 8'h2C;
		16'hCAB7: out_word = 8'hFC;
		16'hCAB8: out_word = 8'h9C;
		16'hCAB9: out_word = 8'h2D;
		16'hCABA: out_word = 8'h6A;
		16'hCABB: out_word = 8'h7D;
		16'hCABC: out_word = 8'h10;
		16'hCABD: out_word = 8'hAF;
		16'hCABE: out_word = 8'hC5;
		16'hCABF: out_word = 8'h3D;
		16'hCAC0: out_word = 8'hD7;
		16'hCAC1: out_word = 8'hEA;
		16'hCAC2: out_word = 8'h1A;
		16'hCAC3: out_word = 8'h92;
		16'hCAC4: out_word = 8'h77;
		16'hCAC5: out_word = 8'hEA;
		16'hCAC6: out_word = 8'hFC;
		16'hCAC7: out_word = 8'hDD;
		16'hCAC8: out_word = 8'hEA;
		16'hCAC9: out_word = 8'h55;
		16'hCACA: out_word = 8'h3E;
		16'hCACB: out_word = 8'h89;
		16'hCACC: out_word = 8'hDF;
		16'hCACD: out_word = 8'hFB;
		16'hCACE: out_word = 8'h1E;
		16'hCACF: out_word = 8'h20;
		16'hCAD0: out_word = 8'h2F;
		16'hCAD1: out_word = 8'h76;
		16'hCAD2: out_word = 8'hED;
		16'hCAD3: out_word = 8'h50;
		16'hCAD4: out_word = 8'h1B;
		16'hCAD5: out_word = 8'h78;
		16'hCAD6: out_word = 8'hBA;
		16'hCAD7: out_word = 8'h03;
		16'hCAD8: out_word = 8'h0F;
		16'hCAD9: out_word = 8'h1D;
		16'hCADA: out_word = 8'h34;
		16'hCADB: out_word = 8'hA6;
		16'hCADC: out_word = 8'h05;
		16'hCADD: out_word = 8'hF7;
		16'hCADE: out_word = 8'hD3;
		16'hCADF: out_word = 8'h28;
		16'hCAE0: out_word = 8'h06;
		16'hCAE1: out_word = 8'hB4;
		16'hCAE2: out_word = 8'hCB;
		16'hCAE3: out_word = 8'hCE;
		16'hCAE4: out_word = 8'h8B;
		16'hCAE5: out_word = 8'hC8;
		16'hCAE6: out_word = 8'h8E;
		16'hCAE7: out_word = 8'hD7;
		16'hCAE8: out_word = 8'h37;
		16'hCAE9: out_word = 8'hC9;
		16'hCAEA: out_word = 8'h88;
		16'hCAEB: out_word = 8'h16;
		16'hCAEC: out_word = 8'h88;
		16'hCAED: out_word = 8'hE8;
		16'hCAEE: out_word = 8'hD9;
		16'hCAEF: out_word = 8'h7F;
		16'hCAF0: out_word = 8'hE8;
		16'hCAF1: out_word = 8'h32;
		16'hCAF2: out_word = 8'hD2;
		16'hCAF3: out_word = 8'h63;
		16'hCAF4: out_word = 8'h93;
		16'hCAF5: out_word = 8'h28;
		16'hCAF6: out_word = 8'h14;
		16'hCAF7: out_word = 8'hC2;
		16'hCAF8: out_word = 8'hF2;
		16'hCAF9: out_word = 8'hE9;
		16'hCAFA: out_word = 8'hFE;
		16'hCAFB: out_word = 8'h85;
		16'hCAFC: out_word = 8'h38;
		16'hCAFD: out_word = 8'h01;
		16'hCAFE: out_word = 8'hAF;
		16'hCAFF: out_word = 8'h6F;
		16'hCB00: out_word = 8'h18;
		16'hCB01: out_word = 8'h0A;
		16'hCB02: out_word = 8'h78;
		16'hCB03: out_word = 8'hF9;
		16'hCB04: out_word = 8'h04;
		16'hCB05: out_word = 8'hFE;
		16'hCB06: out_word = 8'hF9;
		16'hCB07: out_word = 8'h98;
		16'hCB08: out_word = 8'h02;
		16'hCB09: out_word = 8'h3E;
		16'hCB0A: out_word = 8'h93;
		16'hCB0B: out_word = 8'h6F;
		16'hCB0C: out_word = 8'hE1;
		16'hCB0D: out_word = 8'hFF;
		16'hCB0E: out_word = 8'h4F;
		16'hCB0F: out_word = 8'hE1;
		16'hCB10: out_word = 8'hD3;
		16'hCB11: out_word = 8'h63;
		16'hCB12: out_word = 8'h92;
		16'hCB13: out_word = 8'h28;
		16'hCB14: out_word = 8'h81;
		16'hCB15: out_word = 8'h16;
		16'hCB16: out_word = 8'h44;
		16'hCB17: out_word = 8'hF4;
		16'hCB18: out_word = 8'hF2;
		16'hCB19: out_word = 8'h0A;
		16'hCB1A: out_word = 8'h64;
		16'hCB1B: out_word = 8'h84;
		16'hCB1C: out_word = 8'hDF;
		16'hCB1D: out_word = 8'h90;
		16'hCB1E: out_word = 8'h67;
		16'hCB1F: out_word = 8'hDF;
		16'hCB20: out_word = 8'h52;
		16'hCB21: out_word = 8'hDF;
		16'hCB22: out_word = 8'hB8;
		16'hCB23: out_word = 8'h82;
		16'hCB24: out_word = 8'hDF;
		16'hCB25: out_word = 8'h13;
		16'hCB26: out_word = 8'h16;
		16'hCB27: out_word = 8'hBA;
		16'hCB28: out_word = 8'hC9;
		16'hCB29: out_word = 8'hE2;
		16'hCB2A: out_word = 8'hDD;
		16'hCB2B: out_word = 8'h66;
		16'hCB2C: out_word = 8'h01;
		16'hCB2D: out_word = 8'hF9;
		16'hCB2E: out_word = 8'h6E;
		16'hCB2F: out_word = 8'h00;
		16'hCB30: out_word = 8'hED;
		16'hCB31: out_word = 8'h5B;
		16'hCB32: out_word = 8'hF5;
		16'hCB33: out_word = 8'hF1;
		16'hCB34: out_word = 8'h06;
		16'hCB35: out_word = 8'h03;
		16'hCB36: out_word = 8'hCB;
		16'hCB37: out_word = 8'h3A;
		16'hCB38: out_word = 8'hBF;
		16'hCB39: out_word = 8'h3B;
		16'hCB3A: out_word = 8'h10;
		16'hCB3B: out_word = 8'hFA;
		16'hCB3C: out_word = 8'h7B;
		16'hCB3D: out_word = 8'hBD;
		16'hCB3E: out_word = 8'hD8;
		16'hCB3F: out_word = 8'hFC;
		16'hCB40: out_word = 8'h7D;
		16'hCB41: out_word = 8'hDD;
		16'hCB42: out_word = 8'h86;
		16'hCB43: out_word = 8'h03;
		16'hCB44: out_word = 8'h3D;
		16'hCB45: out_word = 8'hBB;
		16'hCB46: out_word = 8'h1E;
		16'hCB47: out_word = 8'h7A;
		16'hCB48: out_word = 8'h24;
		16'hCB49: out_word = 8'hBC;
		16'hCB4A: out_word = 8'h24;
		16'hCB4B: out_word = 8'h7C;
		16'hCB4C: out_word = 8'hF9;
		16'hCB4D: out_word = 8'hF5;
		16'hCB4E: out_word = 8'h02;
		16'hCB4F: out_word = 8'hD6;
		16'hCB50: out_word = 8'h03;
		16'hCB51: out_word = 8'hBA;
		16'hCB52: out_word = 8'hF4;
		16'hCB53: out_word = 8'hCC;
		16'hCB54: out_word = 8'h94;
		16'hCB55: out_word = 8'h4F;
		16'hCB56: out_word = 8'hD8;
		16'hCB57: out_word = 8'h12;
		16'hCB58: out_word = 8'hFA;
		16'hCB59: out_word = 8'hD2;
		16'hCB5A: out_word = 8'h13;
		16'hCB5B: out_word = 8'h06;
		16'hCB5C: out_word = 8'h00;
		16'hCB5D: out_word = 8'h50;
		16'hCB5E: out_word = 8'hEF;
		16'hCB5F: out_word = 8'hE2;
		16'hCB60: out_word = 8'hED;
		16'hCB61: out_word = 8'h52;
		16'hCB62: out_word = 8'h09;
		16'hCB63: out_word = 8'h0A;
		16'hCB64: out_word = 8'h75;
		16'hCB65: out_word = 8'h70;
		16'hCB66: out_word = 8'hF1;
		16'hCB67: out_word = 8'h74;
		16'hCB68: out_word = 8'h13;
		16'hCB69: out_word = 8'hBF;
		16'hCB6A: out_word = 8'h71;
		16'hCB6B: out_word = 8'h0F;
		16'hCB6C: out_word = 8'hC3;
		16'hCB6D: out_word = 8'hE2;
		16'hCB6E: out_word = 8'h7F;
		16'hCB6F: out_word = 8'h01;
		16'hCB70: out_word = 8'h3E;
		16'hCB71: out_word = 8'h73;
		16'hCB72: out_word = 8'h78;
		16'hCB73: out_word = 8'hCD;
		16'hCB74: out_word = 8'hB1;
		16'hCB75: out_word = 8'h22;
		16'hCB76: out_word = 8'h39;
		16'hCB77: out_word = 8'h19;
		16'hCB78: out_word = 8'hAE;
		16'hCB79: out_word = 8'hE5;
		16'hCB7A: out_word = 8'hF4;
		16'hCB7B: out_word = 8'h2C;
		16'hCB7C: out_word = 8'h3E;
		16'hCB7D: out_word = 8'h06;
		16'hCB7E: out_word = 8'h3C;
		16'hCB7F: out_word = 8'h3B;
		16'hCB80: out_word = 8'hFF;
		16'hCB81: out_word = 8'hFE;
		16'hCB82: out_word = 8'h0C;
		16'hCB83: out_word = 8'h20;
		16'hCB84: out_word = 8'h05;
		16'hCB85: out_word = 8'h3E;
		16'hCB86: out_word = 8'h01;
		16'hCB87: out_word = 8'hAE;
		16'hCB88: out_word = 8'h77;
		16'hCB89: out_word = 8'hF9;
		16'hCB8A: out_word = 8'hAF;
		16'hCB8B: out_word = 8'h32;
		16'hCB8C: out_word = 8'h6D;
		16'hCB8D: out_word = 8'h64;
		16'hCB8E: out_word = 8'h3A;
		16'hCB8F: out_word = 8'hA1;
		16'hCB90: out_word = 8'h3E;
		16'hCB91: out_word = 8'h44;
		16'hCB92: out_word = 8'h2F;
		16'hCB93: out_word = 8'hC6;
		16'hCB94: out_word = 8'h09;
		16'hCB95: out_word = 8'h4F;
		16'hCB96: out_word = 8'hEF;
		16'hCB97: out_word = 8'hFA;
		16'hCB98: out_word = 8'h87;
		16'hCB99: out_word = 8'h01;
		16'hCB9A: out_word = 8'h21;
		16'hCB9B: out_word = 8'h20;
		16'hCB9C: out_word = 8'h65;
		16'hCB9D: out_word = 8'hFC;
		16'hCB9E: out_word = 8'h52;
		16'hCB9F: out_word = 8'h30;
		16'hCBA0: out_word = 8'h33;
		16'hCBA1: out_word = 8'h06;
		16'hCBA2: out_word = 8'hD1;
		16'hCBA3: out_word = 8'hFF;
		16'hCBA4: out_word = 8'hC5;
		16'hCBA5: out_word = 8'h41;
		16'hCBA6: out_word = 8'h4E;
		16'hCBA7: out_word = 8'h23;
		16'hCBA8: out_word = 8'hE5;
		16'hCBA9: out_word = 8'h6E;
		16'hCBAA: out_word = 8'hEB;
		16'hCBAB: out_word = 8'h3E;
		16'hCBAC: out_word = 8'hFE;
		16'hCBAD: out_word = 8'hFF;
		16'hCBAE: out_word = 8'h16;
		16'hCBAF: out_word = 8'h00;
		16'hCBB0: out_word = 8'h37;
		16'hCBB1: out_word = 8'hCB;
		16'hCBB2: out_word = 8'h11;
		16'hCBB3: out_word = 8'h17;
		16'hCBB4: out_word = 8'h2C;
		16'hCBB5: out_word = 8'h23;
		16'hCBB6: out_word = 8'h3F;
		16'hCBB7: out_word = 8'h12;
		16'hCBB8: out_word = 8'h10;
		16'hCBB9: out_word = 8'hF6;
		16'hCBBA: out_word = 8'hA6;
		16'hCBBB: out_word = 8'hFC;
		16'hCBBC: out_word = 8'hB2;
		16'hCBBD: out_word = 8'h77;
		16'hCBBE: out_word = 8'h2C;
		16'hCBBF: out_word = 8'h7E;
		16'hCBC0: out_word = 8'hA1;
		16'hCBC1: out_word = 8'hB3;
		16'hCBC2: out_word = 8'h37;
		16'hCBC3: out_word = 8'h7F;
		16'hCBC4: out_word = 8'hEF;
		16'hCBC5: out_word = 8'hEB;
		16'hCBC6: out_word = 8'hE1;
		16'hCBC7: out_word = 8'hF9;
		16'hCBC8: out_word = 8'h23;
		16'hCBC9: out_word = 8'hC1;
		16'hCBCA: out_word = 8'h10;
		16'hCBCB: out_word = 8'hD9;
		16'hCBCC: out_word = 8'hC9;
		16'hCBCD: out_word = 8'h8D;
		16'hCBCE: out_word = 8'h8B;
		16'hCBCF: out_word = 8'h14;
		16'hCBD0: out_word = 8'h56;
		16'hCBD1: out_word = 8'hF0;
		16'hCBD2: out_word = 8'h15;
		16'hCBD3: out_word = 8'h7A;
		16'hCBD4: out_word = 8'hB3;
		16'hCBD5: out_word = 8'hC8;
		16'hCBD6: out_word = 8'hB1;
		16'hCBD7: out_word = 8'hE5;
		16'hCBD8: out_word = 8'hD5;
		16'hCBD9: out_word = 8'h69;
		16'hCBDA: out_word = 8'hE1;
		16'hCBDB: out_word = 8'h01;
		16'hCBDC: out_word = 8'hCB;
		16'hCBDD: out_word = 8'hBD;
		16'hCBDE: out_word = 8'h3C;
		16'hCBDF: out_word = 8'hFE;
		16'hCBE0: out_word = 8'h3D;
		16'hCBE1: out_word = 8'h73;
		16'hCBE2: out_word = 8'hFE;
		16'hCBE3: out_word = 8'hDD;
		16'hCBE4: out_word = 8'h7E;
		16'hCBE5: out_word = 8'hF3;
		16'hCBE6: out_word = 8'h00;
		16'hCBE7: out_word = 8'h3C;
		16'hCBE8: out_word = 8'h28;
		16'hCBE9: out_word = 8'h23;
		16'hCBEA: out_word = 8'h4B;
		16'hCBEB: out_word = 8'hBE;
		16'hCBEC: out_word = 8'hE4;
		16'hCBED: out_word = 8'h01;
		16'hCBEE: out_word = 8'h38;
		16'hCBEF: out_word = 8'h20;
		16'hCBF0: out_word = 8'hF4;
		16'hCBF1: out_word = 8'h33;
		16'hCBF2: out_word = 8'h4E;
		16'hCBF3: out_word = 8'h04;
		16'hCBF4: out_word = 8'hF9;
		16'hCBF5: out_word = 8'h3D;
		16'hCBF6: out_word = 8'hBD;
		16'hCBF7: out_word = 8'h38;
		16'hCBF8: out_word = 8'h16;
		16'hCBF9: out_word = 8'h7C;
		16'hCBFA: out_word = 8'hF0;
		16'hCBFB: out_word = 8'h85;
		16'hCBFC: out_word = 8'h02;
		16'hCBFD: out_word = 8'h10;
		16'hCBFE: out_word = 8'h21;
		16'hCBFF: out_word = 8'hF0;
		16'hCC00: out_word = 8'hB9;
		16'hCC01: out_word = 8'h33;
		16'hCC02: out_word = 8'hBC;
		16'hCC03: out_word = 8'hCC;
		16'hCC04: out_word = 8'h38;
		16'hCC05: out_word = 8'h06;
		16'hCC06: out_word = 8'hF6;
		16'hCC07: out_word = 8'h05;
		16'hCC08: out_word = 8'hE4;
		16'hCC09: out_word = 8'hC6;
		16'hCC0A: out_word = 8'hC9;
		16'hCC0B: out_word = 8'h11;
		16'hCC0C: out_word = 8'h40;
		16'hCC0D: out_word = 8'h2F;
		16'hCC0E: out_word = 8'h19;
		16'hCC0F: out_word = 8'h18;
		16'hCC10: out_word = 8'hCD;
		16'hCC11: out_word = 8'h01;
		16'hCC12: out_word = 8'hFF;
		16'hCC13: out_word = 8'h02;
		16'hCC14: out_word = 8'h03;
		16'hCC15: out_word = 8'h04;
		16'hCC16: out_word = 8'h05;
		16'hCC17: out_word = 8'h06;
		16'hCC18: out_word = 8'h07;
		16'hCC19: out_word = 8'h08;
		16'hCC1A: out_word = 8'h09;
		16'hCC1B: out_word = 8'hFF;
		16'hCC1C: out_word = 8'h0A;
		16'hCC1D: out_word = 8'h0B;
		16'hCC1E: out_word = 8'h0C;
		16'hCC1F: out_word = 8'h0D;
		16'hCC20: out_word = 8'h0E;
		16'hCC21: out_word = 8'h0F;
		16'hCC22: out_word = 8'h10;
		16'hCC23: out_word = 8'h01;
		16'hCC24: out_word = 8'hF0;
		16'hCC25: out_word = 8'h3F;
		16'hCC26: out_word = 8'h00;
		16'hCC27: out_word = 8'h1F;
		16'hCC28: out_word = 8'h40;
		16'hCC29: out_word = 8'h7F;
		16'hCC2A: out_word = 8'h60;
		16'hCC2B: out_word = 8'h07;
		16'hCC2C: out_word = 8'h50;
		16'hCC2D: out_word = 8'h03;
		16'hCC2E: out_word = 8'h48;
		16'hCC2F: out_word = 8'h01;
		16'hCC30: out_word = 8'h8D;
		16'hCC31: out_word = 8'h4C;
		16'hCC32: out_word = 8'h70;
		16'hCC33: out_word = 8'h02;
		16'hCC34: out_word = 8'h00;
		16'hCC35: out_word = 8'hD5;
		16'hCC36: out_word = 8'hF0;
		16'hCC37: out_word = 8'h70;
		16'hCC38: out_word = 8'hF7;
		16'hCC39: out_word = 8'h03;
		16'hCC3A: out_word = 8'h78;
		16'hCC3B: out_word = 8'h01;
		16'hCC3C: out_word = 8'h7C;
		16'hCC3D: out_word = 8'h23;
		16'hCC3E: out_word = 8'hF0;
		16'hCC3F: out_word = 8'h08;
		16'hCC40: out_word = 8'hCF;
		16'hCC41: out_word = 8'h05;
		16'hCC42: out_word = 8'h61;
		16'hCC43: out_word = 8'h3A;
		16'hCC44: out_word = 8'h99;
		16'hCC45: out_word = 8'h65;
		16'hCC46: out_word = 8'hD2;
		16'hCC47: out_word = 8'h20;
		16'hCC48: out_word = 8'h00;
		16'hCC49: out_word = 8'hFF;
		16'hCC4A: out_word = 8'h56;
		16'hCC4B: out_word = 8'h08;
		16'hCC4C: out_word = 8'h50;
		16'hCC4D: out_word = 8'h03;
		16'hCC4E: out_word = 8'h1C;
		16'hCC4F: out_word = 8'hFF;
		16'hCC50: out_word = 8'hFF;
		16'hCC51: out_word = 8'h14;
		16'hCC52: out_word = 8'h01;
		16'hCC53: out_word = 8'h44;
		16'hCC54: out_word = 8'h4F;
		16'hCC55: out_word = 8'h53;
		16'hCC56: out_word = 8'h20;
		16'hCC57: out_word = 8'h4D;
		16'hCC58: out_word = 8'h45;
		16'hCC59: out_word = 8'h0B;
		16'hCC5A: out_word = 8'h49;
		16'hCC5B: out_word = 8'h54;
		16'hCC5C: out_word = 8'h8C;
		16'hCC5D: out_word = 8'h41;
		16'hCC5E: out_word = 8'h17;
		16'hCC5F: out_word = 8'h21;
		16'hCC60: out_word = 8'h14;
		16'hCC61: out_word = 8'h00;
		16'hCC62: out_word = 8'hF1;
		16'hCC63: out_word = 8'h0D;
		16'hCC64: out_word = 8'h20;
		16'hCC65: out_word = 8'h52;
		16'hCC66: out_word = 8'h2E;
		16'hCC67: out_word = 8'hBF;
		16'hCC68: out_word = 8'h65;
		16'hCC69: out_word = 8'h74;
		16'hCC6A: out_word = 8'h72;
		16'hCC6B: out_word = 8'h79;
		16'hCC6C: out_word = 8'h3A;
		16'hCC6D: out_word = 8'h20;
		16'hCC6E: out_word = 8'h4B;
		16'hCC6F: out_word = 8'hFF;
		16'hCC70: out_word = 8'h2F;
		16'hCC71: out_word = 8'h87;
		16'hCC72: out_word = 8'hFD;
		16'hCC73: out_word = 8'hED;
		16'hCC74: out_word = 8'h49;
		16'hCC75: out_word = 8'h2E;
		16'hCC76: out_word = 8'h1B;
		16'hCC77: out_word = 8'h67;
		16'hCC78: out_word = 8'h6E;
		16'hCC79: out_word = 8'hCC;
		16'hCC7A: out_word = 8'h6F;
		16'hCC7B: out_word = 8'h72;
		16'hCC7C: out_word = 8'hC4;
		16'hCC7D: out_word = 8'h73;
		16'hCC7E: out_word = 8'h5C;
		16'hCC7F: out_word = 8'h63;
		16'hCC80: out_word = 8'h74;
		16'hCC81: out_word = 8'h9C;
		16'hCC82: out_word = 8'hF8;
		16'hCC83: out_word = 8'hEF;
		16'hCC84: out_word = 8'h42;
		16'hCC85: out_word = 8'h2E;
		16'hCC86: out_word = 8'h63;
		16'hCC87: out_word = 8'hF2;
		16'hCC88: out_word = 8'h61;
		16'hCC89: out_word = 8'h90;
		16'hCC8A: out_word = 8'h6B;
		16'hCC8B: out_word = 8'hBB;
		16'hCC8C: out_word = 8'hBE;
		16'hCC8D: out_word = 8'h69;
		16'hCC8E: out_word = 8'h62;
		16'hCC8F: out_word = 8'h53;
		16'hCC90: out_word = 8'h86;
		16'hCC91: out_word = 8'h57;
		16'hCC92: out_word = 8'h37;
		16'hCC93: out_word = 8'hF0;
		16'hCC94: out_word = 8'h75;
		16'hCC95: out_word = 8'h08;
		16'hCC96: out_word = 8'h8F;
		16'hCC97: out_word = 8'h0A;
		16'hCC98: out_word = 8'h12;
		16'hCC99: out_word = 8'hF7;
		16'hCC9A: out_word = 8'h0F;
		16'hCC9B: out_word = 8'h1F;
		16'hCC9C: out_word = 8'h6E;
		16'hCC9D: out_word = 8'h66;
		16'hCC9E: out_word = 8'hB2;
		16'hCC9F: out_word = 8'hA1;
		16'hCCA0: out_word = 8'hB5;
		16'hCCA1: out_word = 8'h65;
		16'hCCA2: out_word = 8'h91;
		16'hCCA3: out_word = 8'hD5;
		16'hCCA4: out_word = 8'hA1;
		16'hCCA5: out_word = 8'h53;
		16'hCCA6: out_word = 8'hF8;
		16'hCCA7: out_word = 8'h65;
		16'hCCA8: out_word = 8'h72;
		16'hCCA9: out_word = 8'h76;
		16'hCCAA: out_word = 8'h69;
		16'hCCAB: out_word = 8'h63;
		16'hCCAC: out_word = 8'h76;
		16'hCCAD: out_word = 8'h73;
		16'hCCAE: out_word = 8'hC9;
		16'hCCAF: out_word = 8'hA6;
		16'hCCB0: out_word = 8'h73;
		16'hCCB1: out_word = 8'hA4;
		16'hCCB2: out_word = 8'h02;
		16'hCCB3: out_word = 8'h4E;
		16'hCCB4: out_word = 8'h17;
		16'hCCB5: out_word = 8'h6F;
		16'hCCB6: out_word = 8'h47;
		16'hCCB7: out_word = 8'h53;
		16'hCCB8: out_word = 8'h36;
		16'hCCB9: out_word = 8'hF1;
		16'hCCBA: out_word = 8'h50;
		16'hCCBB: out_word = 8'hAE;
		16'hCCBC: out_word = 8'hF1;
		16'hCCBD: out_word = 8'h70;
		16'hCCBE: out_word = 8'h61;
		16'hCCBF: out_word = 8'h67;
		16'hCCC0: out_word = 8'h42;
		16'hCCC1: out_word = 8'hF8;
		16'hCCC2: out_word = 8'hF3;
		16'hCCC3: out_word = 8'h31;
		16'hCCC4: out_word = 8'h32;
		16'hCCC5: out_word = 8'h38;
		16'hCCC6: out_word = 8'h4B;
		16'hCCC7: out_word = 8'hEC;
		16'hCCC8: out_word = 8'h47;
		16'hCCC9: out_word = 8'h6A;
		16'hCCCA: out_word = 8'hEC;
		16'hCCCB: out_word = 8'hC7;
		16'hCCCC: out_word = 8'h61;
		16'hCCCD: out_word = 8'h6C;
		16'hCCCE: out_word = 8'h68;
		16'hCCCF: out_word = 8'hE8;
		16'hCCD0: out_word = 8'h3D;
		16'hCCD1: out_word = 8'hED;
		16'hCCD2: out_word = 8'h53;
		16'hCCD3: out_word = 8'h2E;
		16'hCCD4: out_word = 8'h43;
		16'hCCD5: out_word = 8'h24;
		16'hCCD6: out_word = 8'h94;
		16'hCCD7: out_word = 8'h74;
		16'hCCD8: out_word = 8'h83;
		16'hCCD9: out_word = 8'h20;
		16'hCCDA: out_word = 8'hFE;
		16'hCCDB: out_word = 8'h6D;
		16'hCCDC: out_word = 8'h64;
		16'hCCDD: out_word = 8'h69;
		16'hCCDE: out_word = 8'h73;
		16'hCCDF: out_word = 8'h6B;
		16'hCCE0: out_word = 8'h04;
		16'hCCE1: out_word = 8'h35;
		16'hCCE2: out_word = 8'h86;
		16'hCCE3: out_word = 8'hD5;
		16'hCCE4: out_word = 8'h6C;
		16'hCCE5: out_word = 8'hE9;
		16'hCCE6: out_word = 8'h4B;
		16'hCCE7: out_word = 8'hE7;
		16'hCCE8: out_word = 8'hE9;
		16'hCCE9: out_word = 8'h36;
		16'hCCEA: out_word = 8'h34;
		16'hCCEB: out_word = 8'h30;
		16'hCCEC: out_word = 8'h4B;
		16'hCCED: out_word = 8'hE9;
		16'hCCEE: out_word = 8'h44;
		16'hCCEF: out_word = 8'h39;
		16'hCCF0: out_word = 8'hE9;
		16'hCCF1: out_word = 8'h37;
		16'hCCF2: out_word = 8'hC3;
		16'hCCF3: out_word = 8'h36;
		16'hCCF4: out_word = 8'h38;
		16'hCCF5: out_word = 8'h46;
		16'hCCF6: out_word = 8'h3E;
		16'hCCF7: out_word = 8'h73;
		16'hCCF8: out_word = 8'hE9;
		16'hCCF9: out_word = 8'h38;
		16'hCCFA: out_word = 8'h39;
		16'hCCFB: out_word = 8'hA4;
		16'hCCFC: out_word = 8'h36;
		16'hCCFD: out_word = 8'hE9;
		16'hCCFE: out_word = 8'h59;
		16'hCCFF: out_word = 8'hF0;
		16'hCD00: out_word = 8'hE9;
		16'hCD01: out_word = 8'h6F;
		16'hCD02: out_word = 8'h70;
		16'hCD03: out_word = 8'h79;
		16'hCD04: out_word = 8'h5C;
		16'hCD05: out_word = 8'hEE;
		16'hCD06: out_word = 8'h23;
		16'hCD07: out_word = 8'h8B;
		16'hCD08: out_word = 8'hA7;
		16'hCD09: out_word = 8'h4A;
		16'hCD0A: out_word = 8'h72;
		16'hCD0B: out_word = 8'h70;
		16'hCD0C: out_word = 8'h67;
		16'hCD0D: out_word = 8'h27;
		16'hCD0E: out_word = 8'hF5;
		16'hCD0F: out_word = 8'hF1;
		16'hCD10: out_word = 8'h79;
		16'hCD11: out_word = 8'hD6;
		16'hCD12: out_word = 8'hF1;
		16'hCD13: out_word = 8'h75;
		16'hCD14: out_word = 8'h48;
		16'hCD15: out_word = 8'h76;
		16'hCD16: out_word = 8'h3F;
		16'hCD17: out_word = 8'hA1;
		16'hCD18: out_word = 8'hA2;
		16'hCD19: out_word = 8'h40;
		16'hCD1A: out_word = 8'hA7;
		16'hCD1B: out_word = 8'h89;
		16'hCD1C: out_word = 8'hAC;
		16'hCD1D: out_word = 8'hB1;
		16'hCD1E: out_word = 8'h0B;
		16'hCD1F: out_word = 8'h10;
		16'hCD20: out_word = 8'h77;
		16'hCD21: out_word = 8'hC9;
		16'hCD22: out_word = 8'h0C;
		16'hCD23: out_word = 8'h05;
		16'hCD24: out_word = 8'h34;
		16'hCD25: out_word = 8'h21;
		16'hCD26: out_word = 8'h2F;
		16'hCD27: out_word = 8'h2F;
		16'hCD28: out_word = 8'h65;
		16'hCD29: out_word = 8'h21;
		16'hCD2A: out_word = 8'h59;
		16'hCD2B: out_word = 8'h9A;
		16'hCD2C: out_word = 8'hFC;
		16'hCD2D: out_word = 8'hBA;
		16'hCD2E: out_word = 8'h21;
		16'hCD2F: out_word = 8'h6C;
		16'hCD30: out_word = 8'hBF;
		16'hCD31: out_word = 8'hED;
		16'hCD32: out_word = 8'h20;
		16'hCD33: out_word = 8'hE6;
		16'hCD34: out_word = 8'h46;
		16'hCD35: out_word = 8'h41;
		16'hCD36: out_word = 8'h54;
		16'hCD37: out_word = 8'hBB;
		16'hCD38: out_word = 8'h65;
		16'hCD39: out_word = 8'hE1;
		16'hCD3A: out_word = 8'h17;
		16'hCD3B: out_word = 8'h18;
		16'hCD3C: out_word = 8'hF3;
		16'hCD3D: out_word = 8'h0F;
		16'hCD3E: out_word = 8'h06;
		16'hCD3F: out_word = 8'h0B;
		16'hCD40: out_word = 8'h0C;
		16'hCD41: out_word = 8'hD5;
		16'hCD42: out_word = 8'h4E;
		16'hCD43: out_word = 8'hBD;
		16'hCD44: out_word = 8'h67;
		16'hCD45: out_word = 8'hD5;
		16'hCD46: out_word = 8'hBF;
		16'hCD47: out_word = 8'h85;
		16'hCD48: out_word = 8'h66;
		16'hCD49: out_word = 8'h09;
		16'hCD4A: out_word = 8'h4C;
		16'hCD4B: out_word = 8'hF9;
		16'hCD4C: out_word = 8'hC0;
		16'hCD4D: out_word = 8'h6A;
		16'hCD4E: out_word = 8'hFF;
		16'hCD4F: out_word = 8'hD5;
		16'hCD50: out_word = 8'h4D;
		16'hCD51: out_word = 8'h61;
		16'hCD52: out_word = 8'h69;
		16'hCD53: out_word = 8'h6E;
		16'hCD54: out_word = 8'h20;
		16'hCD55: out_word = 8'h6D;
		16'hCD56: out_word = 8'h65;
		16'hCD57: out_word = 8'h12;
		16'hCD58: out_word = 8'h75;
		16'hCD59: out_word = 8'hEF;
		16'hCD5A: out_word = 8'hFD;
		16'hCD5B: out_word = 8'hF5;
		16'hCD5C: out_word = 8'h5A;
		16'hCD5D: out_word = 8'h2E;
		16'hCD5E: out_word = 8'h54;
		16'hCD5F: out_word = 8'h52;
		16'hCD60: out_word = 8'h2D;
		16'hCD61: out_word = 8'hDF;
		16'hCD62: out_word = 8'h85;
		16'hCD63: out_word = 8'hC7;
		16'hCD64: out_word = 8'h62;
		16'hCD65: out_word = 8'h6F;
		16'hCD66: out_word = 8'hCD;
		16'hCD67: out_word = 8'h74;
		16'hCD68: out_word = 8'h0D;
		16'hCD69: out_word = 8'hC0;
		16'hCD6A: out_word = 8'h2E;
		16'hCD6B: out_word = 8'h1A;
		16'hCD6C: out_word = 8'hBE;
		16'hCD6D: out_word = 8'h80;
		16'hCD6E: out_word = 8'hF4;
		16'hCD6F: out_word = 8'h39;
		16'hCD70: out_word = 8'hE5;
		16'hCD71: out_word = 8'h61;
		16'hCD72: out_word = 8'h70;
		16'hCD73: out_word = 8'h57;
		16'hCD74: out_word = 8'hC2;
		16'hCD75: out_word = 8'h6C;
		16'hCD76: out_word = 8'h6F;
		16'hCD77: out_word = 8'hBB;
		16'hCD78: out_word = 8'h64;
		16'hCD79: out_word = 8'hF8;
		16'hCD7A: out_word = 8'h97;
		16'hCD7B: out_word = 8'h48;
		16'hCD7C: out_word = 8'h44;
		16'hCD7D: out_word = 8'hEF;
		16'hCD7E: out_word = 8'h3C;
		16'hCD7F: out_word = 8'hE7;
		16'hCD80: out_word = 8'h25;
		16'hCD81: out_word = 8'hD9;
		16'hCD82: out_word = 8'hF5;
		16'hCD83: out_word = 8'h53;
		16'hCD84: out_word = 8'h6A;
		16'hCD85: out_word = 8'hC1;
		16'hCD86: out_word = 8'h72;
		16'hCD87: out_word = 8'h27;
		16'hCD88: out_word = 8'h34;
		16'hCD89: out_word = 8'h4E;
		16'hCD8A: out_word = 8'h20;
		16'hCD8B: out_word = 8'hEA;
		16'hCD8C: out_word = 8'h61;
		16'hCD8D: out_word = 8'h73;
		16'hCD8E: out_word = 8'h4E;
		16'hCD8F: out_word = 8'h84;
		16'hCD90: out_word = 8'hF3;
		16'hCD91: out_word = 8'h55;
		16'hCD92: out_word = 8'h2E;
		16'hCD93: out_word = 8'hBF;
		16'hCD94: out_word = 8'hBA;
		16'hCD95: out_word = 8'h6B;
		16'hCD96: out_word = 8'h79;
		16'hCD97: out_word = 8'h9B;
		16'hCD98: out_word = 8'hDF;
		16'hCD99: out_word = 8'h92;
		16'hCD9A: out_word = 8'h6B;
		16'hCD9B: out_word = 8'hFF;
		16'hCD9C: out_word = 8'h84;
		16'hCD9D: out_word = 8'h00;
		16'hCD9E: out_word = 8'h12;
		16'hCD9F: out_word = 8'h7A;
		16'hCDA0: out_word = 8'h66;
		16'hCDA1: out_word = 8'hE7;
		16'hCDA2: out_word = 8'h74;
		16'hCDA3: out_word = 8'h62;
		16'hCDA4: out_word = 8'h64;
		16'hCDA5: out_word = 8'hDE;
		16'hCDA6: out_word = 8'h75;
		16'hCDA7: out_word = 8'h72;
		16'hCDA8: out_word = 8'hCE;
		16'hCDA9: out_word = 8'h77;
		16'hCDAA: out_word = 8'h6D;
		16'hCDAB: out_word = 8'hDF;
		16'hCDAC: out_word = 8'h33;
		16'hCDAD: out_word = 8'h34;
		16'hCDAE: out_word = 8'h7F;
		16'hCDAF: out_word = 8'h04;
		16'hCDB0: out_word = 8'h76;
		16'hCDB1: out_word = 8'hB2;
		16'hCDB2: out_word = 8'h83;
		16'hCDB3: out_word = 8'hC3;
		16'hCDB4: out_word = 8'h98;
		16'hCDB5: out_word = 8'h2E;
		16'hCDB6: out_word = 8'hC0;
		16'hCDB7: out_word = 8'h75;
		16'hCDB8: out_word = 8'h9E;
		16'hCDB9: out_word = 8'hE2;
		16'hCDBA: out_word = 8'hA8;
		16'hCDBB: out_word = 8'h79;
		16'hCDBC: out_word = 8'h28;
		16'hCDBD: out_word = 8'h42;
		16'hCDBE: out_word = 8'h21;
		16'hCDBF: out_word = 8'h81;
		16'hCDC0: out_word = 8'h15;
		16'hCDC1: out_word = 8'h35;
		16'hCDC2: out_word = 8'h0B;
		16'hCDC3: out_word = 8'h27;
		16'hCDC4: out_word = 8'h62;
		16'hCDC5: out_word = 8'hF6;
		16'hCDC6: out_word = 8'hC0;
		16'hCDC7: out_word = 8'h61;
		16'hCDC8: out_word = 8'h81;
		16'hCDC9: out_word = 8'h85;
		16'hCDCA: out_word = 8'h8E;
		16'hCDCB: out_word = 8'hFE;
		16'hCDCC: out_word = 8'h15;
		16'hCDCD: out_word = 8'h62;
		16'hCDCE: out_word = 8'hF4;
		16'hCDCF: out_word = 8'h40;
		16'hCDD0: out_word = 8'hAF;
		16'hCDD1: out_word = 8'hF1;
		16'hCDD2: out_word = 8'hFF;
		16'hCDD3: out_word = 8'h8C;
		16'hCDD4: out_word = 8'h01;
		16'hCDD5: out_word = 8'h54;
		16'hCDD6: out_word = 8'h1E;
		16'hCDD7: out_word = 8'h18;
		16'hCDD8: out_word = 8'h0A;
		16'hCDD9: out_word = 8'hFE;
		16'hCDDA: out_word = 8'h06;
		16'hCDDB: out_word = 8'h01;
		16'hCDDC: out_word = 8'h38;
		16'hCDDD: out_word = 8'h73;
		16'hCDDE: out_word = 8'hF9;
		16'hCDDF: out_word = 8'hCB;
		16'hCDE0: out_word = 8'h5C;
		16'hCDE1: out_word = 8'hFC;
		16'hCDE2: out_word = 8'hB6;
		16'hCDE3: out_word = 8'h10;
		16'hCDE4: out_word = 8'h98;
		16'hCDE5: out_word = 8'hFE;
		16'hCDE6: out_word = 8'hF8;
		16'hCDE7: out_word = 8'hD0;
		16'hCDE8: out_word = 8'h50;
		16'hCDE9: out_word = 8'hCA;
		16'hCDEA: out_word = 8'h20;
		16'hCDEB: out_word = 8'hCC;
		16'hCDEC: out_word = 8'h4A;
		16'hCDED: out_word = 8'hCF;
		16'hCDEE: out_word = 8'hFE;
		16'hCDEF: out_word = 8'h40;
		16'hCDF0: out_word = 8'hEE;
		16'hCDF1: out_word = 8'hD1;
		16'hCDF2: out_word = 8'hA6;
		16'hCDF3: out_word = 8'hF3;
		16'hCDF4: out_word = 8'hFE;
		16'hCDF5: out_word = 8'h1B;
		16'hCDF6: out_word = 8'h92;
		16'hCDF7: out_word = 8'h0F;
		16'hCDF8: out_word = 8'h10;
		16'hCDF9: out_word = 8'h02;
		16'hCDFA: out_word = 8'h00;
		16'hCDFB: out_word = 8'h6A;
		16'hCDFC: out_word = 8'hFF;
		16'hCDFD: out_word = 8'hCC;
		16'hCDFE: out_word = 8'h01;
		16'hCDFF: out_word = 8'h1A;
		16'hCE00: out_word = 8'hFC;
		16'hCE01: out_word = 8'hC3;
		16'hCE02: out_word = 8'h30;
		16'hCE03: out_word = 8'h29;
		16'hCE04: out_word = 8'h58;
		16'hCE05: out_word = 8'hC2;
		16'hCE06: out_word = 8'h21;
		16'hCE07: out_word = 8'h0A;
		16'hCE08: out_word = 8'h5B;
		16'hCE09: out_word = 8'h2C;
		16'hCE0A: out_word = 8'h17;
		16'hCE0B: out_word = 8'h1E;
		16'hCE0C: out_word = 8'h40;
		16'hCE0D: out_word = 8'hE0;
		16'hCE0E: out_word = 8'h50;
		16'hCE0F: out_word = 8'h14;
		16'hCE10: out_word = 8'h18;
		16'hCE11: out_word = 8'hA1;
		16'hCE12: out_word = 8'hF8;
		16'hCE13: out_word = 8'hBB;
		16'hCE14: out_word = 8'hFE;
		16'hCE15: out_word = 8'h63;
		16'hCE16: out_word = 8'hEC;
		16'hCE17: out_word = 8'hFF;
		16'hCE18: out_word = 8'h57;
		16'hCE19: out_word = 8'hFF;
		16'hCE1A: out_word = 8'hFC;
		16'hCE1B: out_word = 8'hFF;
		16'hCE1C: out_word = 8'hF4;
		16'hCE1D: out_word = 8'h09;
		16'hCE1E: out_word = 8'hA8;
		16'hCE1F: out_word = 8'h10;
		16'hCE20: out_word = 8'h4B;
		16'hCE21: out_word = 8'hFC;
		16'hCE22: out_word = 8'hFB;
		16'hCE23: out_word = 8'hC4;
		16'hCE24: out_word = 8'h15;
		16'hCE25: out_word = 8'h53;
		16'hCE26: out_word = 8'h81;
		16'hCE27: out_word = 8'h0F;
		16'hCE28: out_word = 8'hDC;
		16'hCE29: out_word = 8'hFB;
		16'hCE2A: out_word = 8'h52;
		16'hCE2B: out_word = 8'hF6;
		16'hCE2C: out_word = 8'hC7;
		16'hCE2D: out_word = 8'h50;
		16'hCE2E: out_word = 8'h80;
		16'hCE2F: out_word = 8'hC7;
		16'hCE30: out_word = 8'hEF;
		16'hCE31: out_word = 8'h22;
		16'hCE32: out_word = 8'h84;
		16'hCE33: out_word = 8'h0D;
		16'hCE34: out_word = 8'h6D;
		16'hCE35: out_word = 8'h72;
		16'hCE36: out_word = 8'h20;
		16'hCE37: out_word = 8'h89;
		16'hCE38: out_word = 8'hFF;
		16'hCE39: out_word = 8'hD3;
		16'hCE3A: out_word = 8'h80;
		16'hCE3B: out_word = 8'h67;
		16'hCE3C: out_word = 8'h8F;
		16'hCE3D: out_word = 8'hC1;
		16'hCE3E: out_word = 8'hED;
		16'hCE3F: out_word = 8'h0D;
		16'hCE40: out_word = 8'hCE;
		16'hCE41: out_word = 8'h5C;
		16'hCE42: out_word = 8'hFD;
		16'hCE43: out_word = 8'h06;
		16'hCE44: out_word = 8'h08;
		16'hCE45: out_word = 8'h04;
		16'hCE46: out_word = 8'h14;
		16'hCE47: out_word = 8'h0E;
		16'hCE48: out_word = 8'h0F;
		16'hCE49: out_word = 8'hAB;
		16'hCE4A: out_word = 8'hEF;
		16'hCE4B: out_word = 8'h44;
		16'hCE4C: out_word = 8'h68;
		16'hCE4D: out_word = 8'h6A;
		16'hCE4E: out_word = 8'hF7;
		16'hCE4F: out_word = 8'hDB;
		16'hCE50: out_word = 8'h0D;
		16'hCE51: out_word = 8'h03;
		16'hCE52: out_word = 8'hFF;
		16'hCE53: out_word = 8'hA5;
		16'hCE54: out_word = 8'h69;
		16'hCE55: out_word = 8'h6E;
		16'hCE56: out_word = 8'hC9;
		16'hCE57: out_word = 8'h67;
		16'hCE58: out_word = 8'h2E;
		16'hCE59: out_word = 8'hFF;
		16'hCE5A: out_word = 8'hEF;
		16'hCE5B: out_word = 8'hF1;
		16'hCE5C: out_word = 8'h50;
		16'hCE5D: out_word = 8'h72;
		16'hCE5E: out_word = 8'h65;
		16'hCE5F: out_word = 8'h73;
		16'hCE60: out_word = 8'hE1;
		16'hCE61: out_word = 8'h20;
		16'hCE62: out_word = 8'h70;
		16'hCE63: out_word = 8'h4C;
		16'hCE64: out_word = 8'h41;
		16'hCE65: out_word = 8'h59;
		16'hCE66: out_word = 8'hF0;
		16'hCE67: out_word = 8'h6F;
		16'hCE68: out_word = 8'h6E;
		16'hCE69: out_word = 8'h29;
		16'hCE6A: out_word = 8'h74;
		16'hCE6B: out_word = 8'hE1;
		16'hCE6C: out_word = 8'h00;
		16'hCE6D: out_word = 8'hF1;
		16'hCE6E: out_word = 8'h05;
		16'hCE6F: out_word = 8'h08;
		16'hCE70: out_word = 8'h03;
		16'hCE71: out_word = 8'h16;
		16'hCE72: out_word = 8'hED;
		16'hCE73: out_word = 8'h0F;
		16'hCE74: out_word = 8'h8C;
		16'hCE75: out_word = 8'hB3;
		16'hCE76: out_word = 8'h87;
		16'hCE77: out_word = 8'hC4;
		16'hCE78: out_word = 8'h4E;
		16'hCE79: out_word = 8'h6F;
		16'hCE7A: out_word = 8'h74;
		16'hCE7B: out_word = 8'hB4;
		16'hCE7C: out_word = 8'h20;
		16'hCE7D: out_word = 8'hFB;
		16'hCE7E: out_word = 8'h89;
		16'hCE7F: out_word = 8'hFC;
		16'hCE80: out_word = 8'hCF;
		16'hCE81: out_word = 8'hE2;
		16'hCE82: out_word = 8'hEB;
		16'hCE83: out_word = 8'hFF;
		16'hCE84: out_word = 8'h17;
		16'hCE85: out_word = 8'hA8;
		16'hCE86: out_word = 8'h68;
		16'hCE87: out_word = 8'h12;
		16'hCE88: out_word = 8'h65;
		16'hCE89: out_word = 8'hFB;
		16'hCE8A: out_word = 8'hEC;
		16'hCE8B: out_word = 8'h10;
		16'hCE8C: out_word = 8'h85;
		16'hCE8D: out_word = 8'h61;
		16'hCE8E: out_word = 8'h61;
		16'hCE8F: out_word = 8'hFE;
		16'hCE90: out_word = 8'hA2;
		16'hCE91: out_word = 8'hBA;
		16'hCE92: out_word = 8'hEE;
		16'hCE93: out_word = 8'hCD;
		16'hCE94: out_word = 8'h58;
		16'hCE95: out_word = 8'hBA;
		16'hCE96: out_word = 8'h99;
		16'hCE97: out_word = 8'h5A;
		16'hCE98: out_word = 8'hFF;
		16'hCE99: out_word = 8'h33;
		16'hCE9A: out_word = 8'hCE;
		16'hCE9B: out_word = 8'h03;
		16'hCE9C: out_word = 8'hBA;
		16'hCE9D: out_word = 8'h27;
		16'hCE9E: out_word = 8'hDE;
		16'hCE9F: out_word = 8'h3F;
		16'hCEA0: out_word = 8'h69;
		16'hCEA1: out_word = 8'hC3;
		16'hCEA2: out_word = 8'h82;
		16'hCEA3: out_word = 8'h34;
		16'hCEA4: out_word = 8'hC9;
		16'hCEA5: out_word = 8'h48;
		16'hCEA6: out_word = 8'h4C;
		16'hCEA7: out_word = 8'h20;
		16'hCEA8: out_word = 8'h1E;
		16'hCEA9: out_word = 8'h9F;
		16'hCEAA: out_word = 8'h67;
		16'hCEAB: out_word = 8'h73;
		16'hCEAC: out_word = 8'h00;
		16'hCEAD: out_word = 8'h62;
		16'hCEAE: out_word = 8'h60;
		16'hCEAF: out_word = 8'h8F;
		16'hCEB0: out_word = 8'h08;
		16'hCEB1: out_word = 8'h04;
		16'hCEB2: out_word = 8'hDB;
		16'hCEB3: out_word = 8'h10;
		16'hCEB4: out_word = 8'h17;
		16'hCEB5: out_word = 8'hFD;
		16'hCEB6: out_word = 8'h9C;
		16'hCEB7: out_word = 8'h90;
		16'hCEB8: out_word = 8'hDD;
		16'hCEB9: out_word = 8'h77;
		16'hCEBA: out_word = 8'hA9;
		16'hCEBB: out_word = 8'h9F;
		16'hCEBC: out_word = 8'h6E;
		16'hCEBD: out_word = 8'h25;
		16'hCEBE: out_word = 8'h66;
		16'hCEBF: out_word = 8'h12;
		16'hCEC0: out_word = 8'h75;
		16'hCEC1: out_word = 8'h0D;
		16'hCEC2: out_word = 8'h64;
		16'hCEC3: out_word = 8'hB7;
		16'hCEC4: out_word = 8'hF8;
		16'hCEC5: out_word = 8'hEF;
		16'hCEC6: out_word = 8'h61;
		16'hCEC7: out_word = 8'h6E;
		16'hCEC8: out_word = 8'h79;
		16'hCEC9: out_word = 8'h98;
		16'hCECA: out_word = 8'h6B;
		16'hCECB: out_word = 8'h65;
		16'hCECC: out_word = 8'h96;
		16'hCECD: out_word = 8'h00;
		16'hCECE: out_word = 8'h5A;
		16'hCECF: out_word = 8'hCB;
		16'hCED0: out_word = 8'h8C;
		16'hCED1: out_word = 8'hC8;
		16'hCED2: out_word = 8'h7B;
		16'hCED3: out_word = 8'hCB;
		16'hCED4: out_word = 8'h46;
		16'hCED5: out_word = 8'h69;
		16'hCED6: out_word = 8'h6C;
		16'hCED7: out_word = 8'h65;
		16'hCED8: out_word = 8'h18;
		16'hCED9: out_word = 8'h4F;
		16'hCEDA: out_word = 8'hCA;
		16'hCEDB: out_word = 8'h16;
		16'hCEDC: out_word = 8'hDD;
		16'hCEDD: out_word = 8'h17;
		16'hCEDE: out_word = 8'h04;
		16'hCEDF: out_word = 8'h45;
		16'hCEE0: out_word = 8'hED;
		16'hCEE1: out_word = 8'h56;
		16'hCEE2: out_word = 8'h4F;
		16'hCEE3: out_word = 8'h20;
		16'hCEE4: out_word = 8'h3A;
		16'hCEE5: out_word = 8'h33;
		16'hCEE6: out_word = 8'hD7;
		16'hCEE7: out_word = 8'hC0;
		16'hCEE8: out_word = 8'h78;
		16'hCEE9: out_word = 8'h07;
		16'hCEEA: out_word = 8'h30;
		16'hCEEB: out_word = 8'hC8;
		16'hCEEC: out_word = 8'h2E;
		16'hCEED: out_word = 8'h32;
		16'hCEEE: out_word = 8'hFE;
		16'hCEEF: out_word = 8'h39;
		16'hCEF0: out_word = 8'h16;
		16'hCEF1: out_word = 8'h08;
		16'hCEF2: out_word = 8'hE2;
		16'hCEF3: out_word = 8'hFF;
		16'hCEF4: out_word = 8'h06;
		16'hCEF5: out_word = 8'h5A;
		16'hCEF6: out_word = 8'h58;
		16'hCEF7: out_word = 8'h2D;
		16'hCEF8: out_word = 8'h45;
		16'hCEF9: out_word = 8'h76;
		16'hCEFA: out_word = 8'h6F;
		16'hCEFB: out_word = 8'h6C;
		16'hCEFC: out_word = 8'hEB;
		16'hCEFD: out_word = 8'h75;
		16'hCEFE: out_word = 8'h74;
		16'hCEFF: out_word = 8'h69;
		16'hCF00: out_word = 8'hFE;
		16'hCF01: out_word = 8'h89;
		16'hCF02: out_word = 8'h34;
		16'hCF03: out_word = 8'h30;
		16'hCF04: out_word = 8'h39;
		16'hCF05: out_word = 8'h36;
		16'hCF06: out_word = 8'h1E;
		16'hCF07: out_word = 8'h4B;
		16'hCF08: out_word = 8'h62;
		16'hCF09: out_word = 8'h67;
		16'hCF0A: out_word = 8'hE6;
		16'hCF0B: out_word = 8'h10;
		16'hCF0C: out_word = 8'hE6;
		16'hCF0D: out_word = 8'h45;
		16'hCF0E: out_word = 8'h77;
		16'hCF0F: out_word = 8'h3F;
		16'hCF10: out_word = 8'hFF;
		16'hCF11: out_word = 8'h2E;
		16'hCF12: out_word = 8'h6E;
		16'hCF13: out_word = 8'h65;
		16'hCF14: out_word = 8'h64;
		16'hCF15: out_word = 8'h6F;
		16'hCF16: out_word = 8'hC1;
		16'hCF17: out_word = 8'h70;
		16'hCF18: out_word = 8'h63;
		16'hCF19: out_word = 8'h18;
		16'hCF1A: out_word = 8'h39;
		16'hCF1B: out_word = 8'h6D;
		16'hCF1C: out_word = 8'hEC;
		16'hCF1D: out_word = 8'h9E;
		16'hCF1E: out_word = 8'h18;
		16'hCF1F: out_word = 8'hEC;
		16'hCF20: out_word = 8'h05;
		16'hCF21: out_word = 8'h42;
		16'hCF22: out_word = 8'h61;
		16'hCF23: out_word = 8'hB8;
		16'hCF24: out_word = 8'h86;
		16'hCF25: out_word = 8'h7F;
		16'hCF26: out_word = 8'hD7;
		16'hCF27: out_word = 8'h66;
		16'hCF28: out_word = 8'h3A;
		16'hCF29: out_word = 8'h20;
		16'hCF2A: out_word = 8'h17;
		16'hCF2B: out_word = 8'hFF;
		16'hCF2C: out_word = 8'h4E;
		16'hCF2D: out_word = 8'h8D;
		16'hCF2E: out_word = 8'h4F;
		16'hCF2F: out_word = 8'h45;
		16'hCF30: out_word = 8'h05;
		16'hCF31: out_word = 8'h8C;
		16'hCF32: out_word = 8'hA0;
		16'hCF33: out_word = 8'hFF;
		16'hCF34: out_word = 8'h16;
		16'hCF35: out_word = 8'h27;
		16'hCF36: out_word = 8'hCF;
		16'hCF37: out_word = 8'h41;
		16'hCF38: out_word = 8'h56;
		16'hCF39: out_word = 8'h52;
		16'hCF3A: out_word = 8'h06;
		16'hCF3B: out_word = 8'h42;
		16'hCF3C: out_word = 8'hBA;
		16'hCF3D: out_word = 8'hD5;
		16'hCF3E: out_word = 8'hC2;
		16'hCF3F: out_word = 8'h34;
		16'hCF40: out_word = 8'hCF;
		16'hCF41: out_word = 8'hB0;
		16'hCF42: out_word = 8'hB5;
		16'hCF43: out_word = 8'hCF;
		16'hCF44: out_word = 8'h01;
		16'hCF45: out_word = 8'h3F;
		16'hCF46: out_word = 8'h43;
		16'hCF47: out_word = 8'hE3;
		16'hCF48: out_word = 8'h31;
		16'hCF49: out_word = 8'h2F;
		16'hCF4A: out_word = 8'h32;
		16'hCF4B: out_word = 8'h44;
		16'hCF4C: out_word = 8'h33;
		16'hCF4D: out_word = 8'hCE;
		16'hCF4E: out_word = 8'h34;
		16'hCF4F: out_word = 8'h20;
		16'hCF50: out_word = 8'hEE;
		16'hCF51: out_word = 8'h63;
		16'hCF52: out_word = 8'h68;
		16'hCF53: out_word = 8'h65;
		16'hCF54: out_word = 8'hC0;
		16'hCF55: out_word = 8'h73;
		16'hCF56: out_word = 8'h4B;
		16'hCF57: out_word = 8'h93;
		16'hCF58: out_word = 8'hD0;
		16'hCF59: out_word = 8'h58;
		16'hCF5A: out_word = 8'hFE;
		16'hCF5B: out_word = 8'h64;
		16'hCF5C: out_word = 8'h72;
		16'hCF5D: out_word = 8'h69;
		16'hCF5E: out_word = 8'h76;
		16'hCF5F: out_word = 8'h65;
		16'hCF60: out_word = 8'h73;
		16'hCF61: out_word = 8'hD0;
		16'hCF62: out_word = 8'hB8;
		16'hCF63: out_word = 8'h00;
		16'hCF64: out_word = 8'hD8;
		16'hCF65: out_word = 8'h57;
		16'hCF66: out_word = 8'h4E;
		16'hCF67: out_word = 8'hDE;
		16'hCF68: out_word = 8'h54;
		16'hCF69: out_word = 8'h75;
		16'hCF6A: out_word = 8'h72;
		16'hCF6B: out_word = 8'h57;
		16'hCF6C: out_word = 8'hE9;
		16'hCF6D: out_word = 8'hA1;
		16'hCF6E: out_word = 8'hC9;
		16'hCF6F: out_word = 8'h2F;
		16'hCF70: out_word = 8'hC7;
		16'hCF71: out_word = 8'h66;
		16'hCF72: out_word = 8'h9D;
		16'hCF73: out_word = 8'h2C;
		16'hCF74: out_word = 8'hED;
		16'hCF75: out_word = 8'h20;
		16'hCF76: out_word = 8'h4D;
		16'hCF77: out_word = 8'h04;
		16'hCF78: out_word = 8'hEC;
		16'hCF79: out_word = 8'hFA;
		16'hCF7A: out_word = 8'h65;
		16'hCF7B: out_word = 8'h6D;
		16'hCF7C: out_word = 8'h6F;
		16'hCF7D: out_word = 8'h72;
		16'hCF7E: out_word = 8'h79;
		16'hCF7F: out_word = 8'hF6;
		16'hCF80: out_word = 8'h9D;
		16'hCF81: out_word = 8'h63;
		16'hCF82: out_word = 8'h6B;
		16'hCF83: out_word = 8'h75;
		16'hCF84: out_word = 8'h29;
		16'hCF85: out_word = 8'h38;
		16'hCF86: out_word = 8'h2F;
		16'hCF87: out_word = 8'hD7;
		16'hCF88: out_word = 8'h70;
		16'hCF89: out_word = 8'h2E;
		16'hCF8A: out_word = 8'hE2;
		16'hCF8B: out_word = 8'h17;
		16'hCF8C: out_word = 8'hEF;
		16'hCF8D: out_word = 8'hB8;
		16'hCF8E: out_word = 8'h06;
		16'hCF8F: out_word = 8'h01;
		16'hCF90: out_word = 8'h0D;
		16'hCF91: out_word = 8'h99;
		16'hCF92: out_word = 8'h76;
		16'hCF93: out_word = 8'hFA;
		16'hCF94: out_word = 8'h07;
		16'hCF95: out_word = 8'hFA;
		16'hCF96: out_word = 8'h99;
		16'hCF97: out_word = 8'h77;
		16'hCF98: out_word = 8'hFA;
		16'hCF99: out_word = 8'h08;
		16'hCF9A: out_word = 8'hFA;
		16'hCF9B: out_word = 8'hF4;
		16'hCF9C: out_word = 8'h6D;
		16'hCF9D: out_word = 8'hFF;
		16'hCF9E: out_word = 8'h16;
		16'hCF9F: out_word = 8'h30;
		16'hCFA0: out_word = 8'h87;
		16'hCFA1: out_word = 8'h6A;
		16'hCFA2: out_word = 8'hA0;
		16'hCFA3: out_word = 8'h11;
		16'hCFA4: out_word = 8'hC7;
		16'hCFA5: out_word = 8'hA5;
		16'hCFA6: out_word = 8'h05;
		16'hCFA7: out_word = 8'h52;
		16'hCFA8: out_word = 8'hF1;
		16'hCFA9: out_word = 8'h41;
		16'hCFAA: out_word = 8'h00;
		16'hCFAB: out_word = 8'h16;
		16'hCFAC: out_word = 8'h38;
		16'hCFAD: out_word = 8'h5B;
		16'hCFAE: out_word = 8'h22;
		16'hCFAF: out_word = 8'hA3;
		16'hCFB0: out_word = 8'h4D;
		16'hCFB1: out_word = 8'hD1;
		16'hCFB2: out_word = 8'h64;
		16'hCFB3: out_word = 8'hEA;
		16'hCFB4: out_word = 8'hC4;
		16'hCFB5: out_word = 8'hE9;
		16'hCFB6: out_word = 8'hBA;
		16'hCFB7: out_word = 8'h31;
		16'hCFB8: out_word = 8'hE7;
		16'hCFB9: out_word = 8'h40;
		16'hCFBA: out_word = 8'h5B;
		16'hCFBB: out_word = 8'hA8;
		16'hCFBC: out_word = 8'h9E;
		16'hCFBD: out_word = 8'h4C;
		16'hCFBE: out_word = 8'h9E;
		16'hCFBF: out_word = 8'hF2;
		16'hCFC0: out_word = 8'hD0;
		16'hCFC1: out_word = 8'h2F;
		16'hCFC2: out_word = 8'h9D;
		16'hCFC3: out_word = 8'hF8;
		16'hCFC4: out_word = 8'h8F;
		16'hCFC5: out_word = 8'hD0;
		16'hCFC6: out_word = 8'h17;
		16'hCFC7: out_word = 8'h4E;
		16'hCFC8: out_word = 8'h30;
		16'hCFC9: out_word = 8'hF7;
		16'hCFCA: out_word = 8'h3A;
		16'hCFCB: out_word = 8'hB9;
		16'hCFCC: out_word = 8'hFD;
		16'hCFCD: out_word = 8'h16;
		16'hCFCE: out_word = 8'h08;
		16'hCFCF: out_word = 8'hD0;
		16'hCFD0: out_word = 8'hFB;
		16'hCFD1: out_word = 8'hBC;
		16'hCFD2: out_word = 8'h2E;
		16'hCFD3: out_word = 8'hFD;
		16'hCFD4: out_word = 8'h5E;
		16'hCFD5: out_word = 8'hE1;
		16'hCFD6: out_word = 8'hE5;
		16'hCFD7: out_word = 8'hB7;
		16'hCFD8: out_word = 8'h07;
		16'hCFD9: out_word = 8'h16;
		16'hCFDA: out_word = 8'h15;
		16'hCFDB: out_word = 8'hE5;
		16'hCFDC: out_word = 8'hC4;
		16'hCFDD: out_word = 8'hF5;
		16'hCFDE: out_word = 8'hE5;
		16'hCFDF: out_word = 8'hE0;
		16'hCFE0: out_word = 8'h0D;
		16'hCFE1: out_word = 8'h08;
		16'hCFE2: out_word = 8'h03;
		16'hCFE3: out_word = 8'h42;
		16'hCFE4: out_word = 8'h2E;
		16'hCFE5: out_word = 8'hF8;
		16'hCFE6: out_word = 8'h0B;
		16'hCFE7: out_word = 8'h71;
		16'hCFE8: out_word = 8'h61;
		16'hCFE9: out_word = 8'h6F;
		16'hCFEA: out_word = 8'h70;
		16'hCFEB: out_word = 8'h0F;
		16'hCFEC: out_word = 8'hD7;
		16'hCFED: out_word = 8'hB6;
		16'hCFEE: out_word = 8'h0D;
		16'hCFEF: out_word = 8'hA1;
		16'hCFF0: out_word = 8'h60;
		16'hCFF1: out_word = 8'h8D;
		16'hCFF2: out_word = 8'hB7;
		16'hCFF3: out_word = 8'hBC;
		16'hCFF4: out_word = 8'h12;
		16'hCFF5: out_word = 8'hA6;
		16'hCFF6: out_word = 8'h17;
		16'hCFF7: out_word = 8'h8C;
		16'hCFF8: out_word = 8'h61;
		16'hCFF9: out_word = 8'h62;
		16'hCFFA: out_word = 8'h78;
		16'hCFFB: out_word = 8'hF8;
		16'hCFFC: out_word = 8'hD3;
		16'hCFFD: out_word = 8'hF2;
		16'hCFFE: out_word = 8'hA1;
		16'hCFFF: out_word = 8'hF4;
		16'hD000: out_word = 8'h2E;
		16'hD001: out_word = 8'h5A;
		16'hD002: out_word = 8'h9C;
		16'hD003: out_word = 8'h43;
		16'hD004: out_word = 8'h1B;
		16'hD005: out_word = 8'h74;
		16'hD006: out_word = 8'h72;
		16'hD007: out_word = 8'hF8;
		16'hD008: out_word = 8'hCC;
		16'hD009: out_word = 8'h53;
		16'hD00A: out_word = 8'h44;
		16'hD00B: out_word = 8'h43;
		16'hD00C: out_word = 8'h61;
		16'hD00D: out_word = 8'h3D;
		16'hD00E: out_word = 8'h64;
		16'hD00F: out_word = 8'h3A;
		16'hD010: out_word = 8'h2E;
		16'hD011: out_word = 8'hFB;
		16'hD012: out_word = 8'h3F;
		16'hD013: out_word = 8'hB7;
		16'hD014: out_word = 8'h20;
		16'hD015: out_word = 8'h3B;
		16'hD016: out_word = 8'hF0;
		16'hD017: out_word = 8'h92;
		16'hD018: out_word = 8'h5C;
		16'hD019: out_word = 8'h4E;
		16'hD01A: out_word = 8'h6A;
		16'hD01B: out_word = 8'h9F;
		16'hD01C: out_word = 8'h52;
		16'hD01D: out_word = 8'h41;
		16'hD01E: out_word = 8'h53;
		16'hD01F: out_word = 8'h54;
		16'hD020: out_word = 8'h45;
		16'hD021: out_word = 8'h52;
		16'hD022: out_word = 8'h7B;
		16'hD023: out_word = 8'hF0;
		16'hD024: out_word = 8'h53;
		16'hD025: out_word = 8'h6D;
		16'hD026: out_word = 8'hDB;
		16'hD027: out_word = 8'h75;
		16'hD028: out_word = 8'h63;
		16'hD029: out_word = 8'h1B;
		16'hD02A: out_word = 8'hF0;
		16'hD02B: out_word = 8'h8F;
		16'hD02C: out_word = 8'hE0;
		16'hD02D: out_word = 8'hCF;
		16'hD02E: out_word = 8'h4C;
		16'hD02F: out_word = 8'h41;
		16'hD030: out_word = 8'h56;
		16'hD031: out_word = 8'hB7;
		16'hD032: out_word = 8'h45;
		16'hD033: out_word = 8'h36;
		16'hD034: out_word = 8'hE0;
		16'hD035: out_word = 8'h2E;
		16'hD036: out_word = 8'hF0;
		16'hD037: out_word = 8'h17;
		16'hD038: out_word = 8'h04;
		16'hD039: out_word = 8'h3B;
		16'hD03A: out_word = 8'h29;
		16'hD03B: out_word = 8'hFB;
		16'hD03C: out_word = 8'h36;
		16'hD03D: out_word = 8'hFB;
		16'hD03E: out_word = 8'h33;
		16'hD03F: out_word = 8'hEF;
		16'hD040: out_word = 8'h32;
		16'hD041: out_word = 8'h20;
		16'hD042: out_word = 8'h02;
		16'hD043: out_word = 8'hEC;
		16'hD044: out_word = 8'h2A;
		16'hD045: out_word = 8'hAA;
		16'hD046: out_word = 8'h29;
		16'hD047: out_word = 8'h01;
		16'hD048: out_word = 8'h44;
		16'hD049: out_word = 8'hE5;
		16'hD04A: out_word = 8'hF0;
		16'hD04B: out_word = 8'h0D;
		16'hD04C: out_word = 8'h10;
		16'hD04D: out_word = 8'hF6;
		16'hD04E: out_word = 8'h93;
		16'hD04F: out_word = 8'hDF;
		16'hD050: out_word = 8'h10;
		16'hD051: out_word = 8'h52;
		16'hD052: out_word = 8'h41;
		16'hD053: out_word = 8'h4D;
		16'hD054: out_word = 8'h44;
		16'hD055: out_word = 8'hFF;
		16'hD056: out_word = 8'h49;
		16'hD057: out_word = 8'h53;
		16'hD058: out_word = 8'h4B;
		16'hD059: out_word = 8'h20;
		16'hD05A: out_word = 8'h06;
		16'hD05B: out_word = 8'h0C;
		16'hD05C: out_word = 8'h03;
		16'hD05D: out_word = 8'h14;
		16'hD05E: out_word = 8'hF3;
		16'hD05F: out_word = 8'h27;
		16'hD060: out_word = 8'h49;
		16'hD061: out_word = 8'h4E;
		16'hD062: out_word = 8'h53;
		16'hD063: out_word = 8'hA2;
		16'hD064: out_word = 8'h54;
		16'hD065: out_word = 8'hE2;
		16'hD066: out_word = 8'h20;
		16'hD067: out_word = 8'h4F;
		16'hD068: out_word = 8'h55;
		16'hD069: out_word = 8'h45;
		16'hD06A: out_word = 8'h50;
		16'hD06B: out_word = 8'h3F;
		16'hD06C: out_word = 8'hF9;
		16'hD06D: out_word = 8'h31;
		16'hD06E: out_word = 8'h2D;
		16'hD06F: out_word = 8'hB4;
		16'hD070: out_word = 8'hFF;
		16'hD071: out_word = 8'h03;
		16'hD072: out_word = 8'h3E;
		16'hD073: out_word = 8'h2E;
		16'hD074: out_word = 8'h1A;
		16'hD075: out_word = 8'hEA;
		16'hD076: out_word = 8'h47;
		16'hD077: out_word = 8'h4F;
		16'hD078: out_word = 8'h91;
		16'hD079: out_word = 8'hA8;
		16'hD07A: out_word = 8'h45;
		16'hD07B: out_word = 8'hF3;
		16'hD07C: out_word = 8'h50;
		16'hD07D: out_word = 8'h2C;
		16'hD07E: out_word = 8'h83;
		16'hD07F: out_word = 8'h55;
		16'hD080: out_word = 8'h0F;
		16'hD081: out_word = 8'h49;
		16'hD082: out_word = 8'h44;
		16'hD083: out_word = 8'h86;
		16'hD084: out_word = 8'h20;
		16'hD085: out_word = 8'h91;
		16'hD086: out_word = 8'hDA;
		16'hD087: out_word = 8'h21;
		16'hD088: out_word = 8'hFF;
		16'hD089: out_word = 8'hA1;
		16'hD08A: out_word = 8'hFF;
		16'hD08B: out_word = 8'h20;
		16'hD08C: out_word = 8'h62;
		16'hD08D: out_word = 8'h65;
		16'hD08E: out_word = 8'h74;
		16'hD08F: out_word = 8'hAF;
		16'hD090: out_word = 8'h61;
		16'hD091: out_word = 8'hAF;
		16'hD092: out_word = 8'hB9;
		16'hD093: out_word = 8'hAF;
		16'hD094: out_word = 8'hCF;
		16'hD095: out_word = 8'hB5;
		16'hD096: out_word = 8'h65;
		16'hD097: out_word = 8'hE0;
		16'hD098: out_word = 8'h56;
		16'hD099: out_word = 8'h30;
		16'hD09A: out_word = 8'h23;
		16'hD09B: out_word = 8'h3F;
		16'hD09C: out_word = 8'hFD;
		16'hD09D: out_word = 8'hB0;
		16'hD09E: out_word = 8'h22;
		16'hD09F: out_word = 8'h36;
		16'hD0A0: out_word = 8'h35;
		16'hD0A1: out_word = 8'h33;
		16'hD0A2: out_word = 8'h16;
		16'hD0A3: out_word = 8'h38;
		16'hD0A4: out_word = 8'h17;
		16'hD0A5: out_word = 8'h3A;
		16'hD0A6: out_word = 8'hF9;
		16'hD0A7: out_word = 8'hC0;
		16'hD0A8: out_word = 8'h3C;
		16'hD0A9: out_word = 8'hF5;
		16'hD0AA: out_word = 8'h31;
		16'hD0AB: out_word = 8'h35;
		16'hD0AC: out_word = 8'h36;
		16'hD0AD: out_word = 8'h59;
		16'hD0AE: out_word = 8'h39;
		16'hD0AF: out_word = 8'hF5;
		16'hD0B0: out_word = 8'h8D;
		16'hD0B1: out_word = 8'hEA;
		16'hD0B2: out_word = 8'hF7;
		16'hD0B3: out_word = 8'h0D;
		16'hD0B4: out_word = 8'hB7;
		16'hD0B5: out_word = 8'h97;
		16'hD0B6: out_word = 8'h08;
		16'hD0B7: out_word = 8'h2F;
		16'hD0B8: out_word = 8'h8B;
		16'hD0B9: out_word = 8'h10;
		16'hD0BA: out_word = 8'h77;
		16'hD0BB: out_word = 8'hF7;
		16'hD0BC: out_word = 8'h0F;
		16'hD0BD: out_word = 8'h36;
		16'hD0BE: out_word = 8'hF0;
		16'hD0BF: out_word = 8'h2C;
		16'hD0C0: out_word = 8'hCC;
		16'hD0C1: out_word = 8'h09;
		16'hD0C2: out_word = 8'h9E;
		16'hD0C3: out_word = 8'h78;
		16'hD0C4: out_word = 8'h93;
		16'hD0C5: out_word = 8'h40;
		16'hD0C6: out_word = 8'h08;
		16'hD0C7: out_word = 8'h18;
		16'hD0C8: out_word = 8'h60;
		16'hD0C9: out_word = 8'hDF;
		16'hD0CA: out_word = 8'h3C;
		16'hD0CB: out_word = 8'h77;
		16'hD0CC: out_word = 8'hB8;
		16'hD0CD: out_word = 8'h7C;
		16'hD0CE: out_word = 8'h7F;
		16'hD0CF: out_word = 8'h8B;
		16'hD0D0: out_word = 8'hF8;
		16'hD0D1: out_word = 8'hC7;
		16'hD0D2: out_word = 8'h89;
		16'hD0D3: out_word = 8'h8C;
		16'hD0D4: out_word = 8'hE3;
		16'hD0D5: out_word = 8'hF9;
		16'hD0D6: out_word = 8'h1C;
		16'hD0D7: out_word = 8'hF0;
		16'hD0D8: out_word = 8'hFF;
		16'hD0D9: out_word = 8'hFC;
		16'hD0DA: out_word = 8'h70;
		16'hD0DB: out_word = 8'hF4;
		16'hD0DC: out_word = 8'hFE;
		16'hD0DD: out_word = 8'h78;
		16'hD0DE: out_word = 8'h1F;
		16'hD0DF: out_word = 8'hE0;
		16'hD0E0: out_word = 8'h3C;
		16'hD0E1: out_word = 8'h07;
		16'hD0E2: out_word = 8'h80;
		16'hD0E3: out_word = 8'h0E;
		16'hD0E4: out_word = 8'hBA;
		16'hD0E5: out_word = 8'h69;
		16'hD0E6: out_word = 8'hB3;
		16'hD0E7: out_word = 8'h98;
		16'hD0E8: out_word = 8'h83;
		16'hD0E9: out_word = 8'h33;
		16'hD0EA: out_word = 8'hFD;
		16'hD0EB: out_word = 8'h87;
		16'hD0EC: out_word = 8'h2E;
		16'hD0ED: out_word = 8'h47;
		16'hD0EE: out_word = 8'h24;
		16'hD0EF: out_word = 8'hFD;
		16'hD0F0: out_word = 8'hEE;
		16'hD0F1: out_word = 8'h2C;
		16'hD0F2: out_word = 8'h4F;
		16'hD0F3: out_word = 8'hC0;
		16'hD0F4: out_word = 8'h22;
		16'hD0F5: out_word = 8'hE5;
		16'hD0F6: out_word = 8'h84;
		16'hD0F7: out_word = 8'hFD;
		16'hD0F8: out_word = 8'hB4;
		16'hD0F9: out_word = 8'hC9;
		16'hD0FA: out_word = 8'hF7;
		16'hD0FB: out_word = 8'h3F;
		16'hD0FC: out_word = 8'hB2;
		16'hD0FD: out_word = 8'hD6;
		16'hD0FE: out_word = 8'h63;
		16'hD0FF: out_word = 8'hA0;
		16'hD100: out_word = 8'hB8;
		16'hD101: out_word = 8'h18;
		16'hD102: out_word = 8'h5A;
		16'hD103: out_word = 8'hB8;
		16'hD104: out_word = 8'hD9;
		16'hD105: out_word = 8'h80;
		16'hD106: out_word = 8'h04;
		16'hD107: out_word = 8'h6D;
		16'hD108: out_word = 8'hB8;
		16'hD109: out_word = 8'hF3;
		16'hD10A: out_word = 8'h3C;
		16'hD10B: out_word = 8'hA8;
		16'hD10C: out_word = 8'hB8;
		16'hD10D: out_word = 8'hEC;
		16'hD10E: out_word = 8'hEA;
		16'hD10F: out_word = 8'h3C;
		16'hD110: out_word = 8'h04;
		16'hD111: out_word = 8'h2A;
		16'hD112: out_word = 8'h1E;
		16'hD113: out_word = 8'hB8;
		16'hD114: out_word = 8'hFF;
		16'hD115: out_word = 8'h18;
		16'hD116: out_word = 8'hC0;
		16'hD117: out_word = 8'h0C;
		16'hD118: out_word = 8'hD5;
		16'hD119: out_word = 8'hB8;
		16'hD11A: out_word = 8'hC3;
		16'hD11B: out_word = 8'h88;
		16'hD11C: out_word = 8'h0C;
		16'hD11D: out_word = 8'h5C;
		16'hD11E: out_word = 8'hBB;
		16'hD11F: out_word = 8'hB8;
		16'hD120: out_word = 8'h8E;
		16'hD121: out_word = 8'h78;
		16'hD122: out_word = 8'hD4;
		16'hD123: out_word = 8'hB8;
		16'hD124: out_word = 8'h4B;
		16'hD125: out_word = 8'hBB;
		16'hD126: out_word = 8'hFE;
		16'hD127: out_word = 8'h0A;
		16'hD128: out_word = 8'h5F;
		16'hD129: out_word = 8'hB8;
		16'hD12A: out_word = 8'h3D;
		16'hD12B: out_word = 8'hF7;
		16'hD12C: out_word = 8'hBE;
		16'hD12D: out_word = 8'h7C;
		16'hD12E: out_word = 8'h4F;
		16'hD12F: out_word = 8'h8A;
		16'hD130: out_word = 8'hC8;
		16'hD131: out_word = 8'h5C;
		16'hD132: out_word = 8'h73;
		16'hD133: out_word = 8'hB8;
		16'hD134: out_word = 8'hC6;
		16'hD135: out_word = 8'h70;
		16'hD136: out_word = 8'h38;
		16'hD137: out_word = 8'h2E;
		16'hD138: out_word = 8'hBB;
		16'hD139: out_word = 8'h72;
		16'hD13A: out_word = 8'hB8;
		16'hD13B: out_word = 8'h08;
		16'hD13C: out_word = 8'h40;
		16'hD13D: out_word = 8'h0E;
		16'hD13E: out_word = 8'hC7;
		16'hD13F: out_word = 8'hC0;
		16'hD140: out_word = 8'hB8;
		16'hD141: out_word = 8'h31;
		16'hD142: out_word = 8'hB8;
		16'hD143: out_word = 8'hFF;
		16'hD144: out_word = 8'hB0;
		16'hD145: out_word = 8'hE0;
		16'hD146: out_word = 8'hFF;
		16'hD147: out_word = 8'hEC;
		16'hD148: out_word = 8'h50;
		16'hD149: out_word = 8'h1A;
		16'hD14A: out_word = 8'hFC;
		16'hD14B: out_word = 8'hC0;
		16'hD14C: out_word = 8'hEE;
		16'hD14D: out_word = 8'h1C;
		16'hD14E: out_word = 8'h5E;
		16'hD14F: out_word = 8'hFC;
		16'hD150: out_word = 8'h0E;
		16'hD151: out_word = 8'h0D;
		16'hD152: out_word = 8'h7D;
		16'hD153: out_word = 8'h10;
		16'hD154: out_word = 8'h01;
		16'hD155: out_word = 8'hAF;
		16'hD156: out_word = 8'h60;
		16'hD157: out_word = 8'hE6;
		16'hD158: out_word = 8'h06;
		16'hD159: out_word = 8'h4B;
		16'hD15A: out_word = 8'h0B;
		16'hD15B: out_word = 8'hFA;
		16'hD15C: out_word = 8'hD6;
		16'hD15D: out_word = 8'hF8;
		16'hD15E: out_word = 8'h10;
		16'hD15F: out_word = 8'hE5;
		16'hD160: out_word = 8'h0B;
		16'hD161: out_word = 8'h4F;
		16'hD162: out_word = 8'hB9;
		16'hD163: out_word = 8'h3E;
		16'hD164: out_word = 8'h14;
		16'hD165: out_word = 8'hED;
		16'hD166: out_word = 8'h79;
		16'hD167: out_word = 8'hFB;
		16'hD168: out_word = 8'hC3;
		16'hD169: out_word = 8'h00;
		16'hD16A: out_word = 8'hC0;
		16'hD16B: out_word = 8'h18;
		16'hD16C: out_word = 8'hF4;
		16'hD16D: out_word = 8'hD9;
		16'hD16E: out_word = 8'hEF;
		16'hD16F: out_word = 8'h3C;
		16'hD170: out_word = 8'h40;
		16'hD171: out_word = 8'hCA;
		16'hD172: out_word = 8'hF7;
		16'hD173: out_word = 8'hCC;
		16'hD174: out_word = 8'h01;
		16'hD175: out_word = 8'hFC;
		16'hD176: out_word = 8'h5F;
		16'hD177: out_word = 8'h83;
		16'hD178: out_word = 8'hCE;
		16'hD179: out_word = 8'h83;
		16'hD17A: out_word = 8'h28;
		16'hD17B: out_word = 8'h02;
		16'hD17C: out_word = 8'h9C;
		16'hD17D: out_word = 8'h07;
		16'hD17E: out_word = 8'hFA;
		16'hD17F: out_word = 8'hB4;
		16'hD180: out_word = 8'h5D;
		16'hD181: out_word = 8'hC4;
		16'hD182: out_word = 8'hFC;
		16'hD183: out_word = 8'h26;
		16'hD184: out_word = 8'h30;
		16'hD185: out_word = 8'hFE;
		16'hD186: out_word = 8'h3B;
		16'hD187: out_word = 8'h0C;
		16'hD188: out_word = 8'hF6;
		16'hD189: out_word = 8'h3A;
		16'hD18A: out_word = 8'h0A;
		16'hD18B: out_word = 8'hB5;
		16'hD18C: out_word = 8'h52;
		16'hD18D: out_word = 8'hFE;
		16'hD18E: out_word = 8'hB3;
		16'hD18F: out_word = 8'hEE;
		16'hD190: out_word = 8'hB7;
		16'hD191: out_word = 8'h05;
		16'hD192: out_word = 8'hC3;
		16'hD193: out_word = 8'h2C;
		16'hD194: out_word = 8'hFE;
		16'hD195: out_word = 8'h2D;
		16'hD196: out_word = 8'hAC;
		16'hD197: out_word = 8'h70;
		16'hD198: out_word = 8'hD8;
		16'hD199: out_word = 8'hB6;
		16'hD19A: out_word = 8'h1A;
		16'hD19B: out_word = 8'h92;
		16'hD19C: out_word = 8'h20;
		16'hD19D: out_word = 8'h93;
		16'hD19E: out_word = 8'h31;
		16'hD19F: out_word = 8'h1C;
		16'hD1A0: out_word = 8'h12;
		16'hD1A1: out_word = 8'hD8;
		16'hD1A2: out_word = 8'hBB;
		16'hD1A3: out_word = 8'hFE;
		16'hD1A4: out_word = 8'hC7;
		16'hD1A5: out_word = 8'hDB;
		16'hD1A6: out_word = 8'hFF;
		16'hD1A7: out_word = 8'hFF;
		16'hD1A8: out_word = 8'h5F;
		16'hD1A9: out_word = 8'h33;
		16'hD1AA: out_word = 8'h1D;
		16'hD1AB: out_word = 8'hD8;
		16'hD1AC: out_word = 8'hC9;
		16'hD1AD: out_word = 8'hBC;
		16'hD1AE: out_word = 8'h74;
		16'hD1AF: out_word = 8'h28;
		16'hD1B0: out_word = 8'hF6;
		16'hD1B1: out_word = 8'h83;
		16'hD1B2: out_word = 8'hFF;
		16'hD1B3: out_word = 8'h8B;
		16'hD1B4: out_word = 8'hE3;
		16'hD1B5: out_word = 8'hA3;
		16'hD1B6: out_word = 8'h3A;
		16'hD1B7: out_word = 8'h39;
		16'hD1B8: out_word = 8'h09;
		16'hD1B9: out_word = 8'h6B;
		16'hD1BA: out_word = 8'hC6;
		16'hD1BB: out_word = 8'h5E;
		16'hD1BC: out_word = 8'h95;
		16'hD1BD: out_word = 8'h07;
		16'hD1BE: out_word = 8'h25;
		16'hD1BF: out_word = 8'h73;
		16'hD1C0: out_word = 8'h8D;
		16'hD1C1: out_word = 8'h74;
		16'hD1C2: out_word = 8'h35;
		16'hD1C3: out_word = 8'hFE;
		16'hD1C4: out_word = 8'h2E;
		16'hD1C5: out_word = 8'h31;
		16'hD1C6: out_word = 8'h61;
		16'hD1C7: out_word = 8'h20;
		16'hD1C8: out_word = 8'h43;
		16'hD1C9: out_word = 8'h00;
		16'hD1CA: out_word = 8'hDB;
		16'hD1CB: out_word = 8'h47;
		16'hD1CC: out_word = 8'hF3;
		16'hD1CD: out_word = 8'hB6;
		16'hD1CE: out_word = 8'h03;
		16'hD1CF: out_word = 8'hE8;
		16'hD1D0: out_word = 8'h3F;
		16'hD1D1: out_word = 8'h17;
		16'hD1D2: out_word = 8'h0B;
		16'hD1D3: out_word = 8'h29;
		16'hD1D4: out_word = 8'hFA;
		16'hD1D5: out_word = 8'h08;
		16'hD1D6: out_word = 8'hFF;
		16'hD1D7: out_word = 8'h80;
		16'hD1D8: out_word = 8'h0F;
		16'hD1D9: out_word = 8'h25;
		16'hD1DA: out_word = 8'h5D;
		16'hD1DB: out_word = 8'hA3;
		16'hD1DC: out_word = 8'h94;
		16'hD1DD: out_word = 8'h5B;
		16'hD1DE: out_word = 8'h43;
		16'hD1DF: out_word = 8'hE6;
		16'hD1E0: out_word = 8'hFF;
		16'hD1E1: out_word = 8'hF4;
		16'hD1E2: out_word = 8'h89;
		16'hD1E3: out_word = 8'h90;
		16'hD1E4: out_word = 8'h5D;
		16'hD1E5: out_word = 8'h2A;
		16'hD1E6: out_word = 8'hF4;
		16'hD1E7: out_word = 8'h2C;
		16'hD1E8: out_word = 8'hAA;
		16'hD1E9: out_word = 8'h28;
		16'hD1EA: out_word = 8'hF0;
		16'hD1EB: out_word = 8'h02;
		16'hD1EC: out_word = 8'hE6;
		16'hD1ED: out_word = 8'h5F;
		16'hD1EE: out_word = 8'h03;
		16'hD1EF: out_word = 8'h6B;
		16'hD1F0: out_word = 8'hFE;
		16'hD1F1: out_word = 8'h01;
		16'hD1F2: out_word = 8'h86;
		16'hD1F3: out_word = 8'hB1;
		16'hD1F4: out_word = 8'h4C;
		16'hD1F5: out_word = 8'h18;
		16'hD1F6: out_word = 8'h68;
		16'hD1F7: out_word = 8'hDE;
		16'hD1F8: out_word = 8'h30;
		16'hD1F9: out_word = 8'hBF;
		16'hD1FA: out_word = 8'hE7;
		16'hD1FB: out_word = 8'hC3;
		16'hD1FC: out_word = 8'hA7;
		16'hD1FD: out_word = 8'h3A;
		16'hD1FE: out_word = 8'hD9;
		16'hD1FF: out_word = 8'h4A;
		16'hD200: out_word = 8'hFC;
		16'hD201: out_word = 8'hDA;
		16'hD202: out_word = 8'h2E;
		16'hD203: out_word = 8'hFC;
		16'hD204: out_word = 8'h78;
		16'hD205: out_word = 8'hAF;
		16'hD206: out_word = 8'h32;
		16'hD207: out_word = 8'h34;
		16'hD208: out_word = 8'h35;
		16'hD209: out_word = 8'h37;
		16'hD20A: out_word = 8'hCF;
		16'hD20B: out_word = 8'hE1;
		16'hD20C: out_word = 8'hAF;
		16'hD20D: out_word = 8'hF5;
		16'hD20E: out_word = 8'hE9;
		16'hD20F: out_word = 8'h33;
		16'hD210: out_word = 8'h39;
		16'hD211: out_word = 8'h30;
		16'hD212: out_word = 8'hF5;
		16'hD213: out_word = 8'hEA;
		16'hD214: out_word = 8'hFE;
		16'hD215: out_word = 8'hED;
		16'hD216: out_word = 8'h5B;
		16'hD217: out_word = 8'hF4;
		16'hD218: out_word = 8'h5C;
		16'hD219: out_word = 8'h01;
		16'hD21A: out_word = 8'h05;
		16'hD21B: out_word = 8'h2E;
		16'hD21C: out_word = 8'h7F;
		16'hD21D: out_word = 8'h17;
		16'hD21E: out_word = 8'h60;
		16'hD21F: out_word = 8'hE5;
		16'hD220: out_word = 8'hC3;
		16'hD221: out_word = 8'h13;
		16'hD222: out_word = 8'h3D;
		16'hD223: out_word = 8'h0D;
		16'hD224: out_word = 8'hFF;
		16'hD225: out_word = 8'hF3;
		16'hD226: out_word = 8'hA7;
		16'hD227: out_word = 8'h21;
		16'hD228: out_word = 8'h4B;
		16'hD229: out_word = 8'h45;
		16'hD22A: out_word = 8'h28;
		16'hD22B: out_word = 8'h0F;
		16'hD22C: out_word = 8'h3D;
		16'hD22D: out_word = 8'h0A;
		16'hD22E: out_word = 8'hF2;
		16'hD22F: out_word = 8'h67;
		16'hD230: out_word = 8'hFA;
		16'hD231: out_word = 8'h09;
		16'hD232: out_word = 8'hFA;
		16'hD233: out_word = 8'h5A;
		16'hD234: out_word = 8'h46;
		16'hD235: out_word = 8'h54;
		16'hD236: out_word = 8'hAE;
		16'hD237: out_word = 8'h87;
		16'hD238: out_word = 8'hC9;
		16'hD239: out_word = 8'h22;
		16'hD23A: out_word = 8'hFF;
		16'hD23B: out_word = 8'hFA;
		16'hD23C: out_word = 8'h43;
		16'hD23D: out_word = 8'h08;
		16'hD23E: out_word = 8'hA7;
		16'hD23F: out_word = 8'h3E;
		16'hD240: out_word = 8'hE0;
		16'hD241: out_word = 8'h28;
		16'hD242: out_word = 8'h02;
		16'hD243: out_word = 8'h13;
		16'hD244: out_word = 8'hF0;
		16'hD245: out_word = 8'h32;
		16'hD246: out_word = 8'hCF;
		16'hD247: out_word = 8'h64;
		16'hD248: out_word = 8'h46;
		16'hD249: out_word = 8'hBA;
		16'hD24A: out_word = 8'h47;
		16'hD24B: out_word = 8'hCD;
		16'hD24C: out_word = 8'hBA;
		16'hD24D: out_word = 8'h8B;
		16'hD24E: out_word = 8'h44;
		16'hD24F: out_word = 8'h40;
		16'hD250: out_word = 8'hF0;
		16'hD251: out_word = 8'h45;
		16'hD252: out_word = 8'hD9;
		16'hD253: out_word = 8'h2A;
		16'hD254: out_word = 8'h09;
		16'hD255: out_word = 8'hF8;
		16'hD256: out_word = 8'h22;
		16'hD257: out_word = 8'hC8;
		16'hD258: out_word = 8'h43;
		16'hD259: out_word = 8'h53;
		16'hD25A: out_word = 8'h0B;
		16'hD25B: out_word = 8'hFA;
		16'hD25C: out_word = 8'hAD;
		16'hD25D: out_word = 8'h0A;
		16'hD25E: out_word = 8'h11;
		16'hD25F: out_word = 8'h3F;
		16'hD260: out_word = 8'h00;
		16'hD261: out_word = 8'h19;
		16'hD262: out_word = 8'h7D;
		16'hD263: out_word = 8'hFF;
		16'hD264: out_word = 8'hA7;
		16'hD265: out_word = 8'h28;
		16'hD266: out_word = 8'h01;
		16'hD267: out_word = 8'h24;
		16'hD268: out_word = 8'h7C;
		16'hD269: out_word = 8'hCB;
		16'hD26A: out_word = 8'h3F;
		16'hD26B: out_word = 8'hCE;
		16'hD26C: out_word = 8'hF1;
		16'hD26D: out_word = 8'h00;
		16'hD26E: out_word = 8'h3D;
		16'hD26F: out_word = 8'hD9;
		16'hD270: out_word = 8'hCA;
		16'hD271: out_word = 8'hF8;
		16'hD272: out_word = 8'h43;
		16'hD273: out_word = 8'hDD;
		16'hD274: out_word = 8'h6F;
		16'hD275: out_word = 8'h58;
		16'hD276: out_word = 8'hCD;
		16'hD277: out_word = 8'hEC;
		16'hD278: out_word = 8'h50;
		16'hD279: out_word = 8'hD5;
		16'hD27A: out_word = 8'hF3;
		16'hD27B: out_word = 8'h21;
		16'hD27C: out_word = 8'h01;
		16'hD27D: out_word = 8'hE5;
		16'hD27E: out_word = 8'hEB;
		16'hD27F: out_word = 8'h87;
		16'hD280: out_word = 8'h30;
		16'hD281: out_word = 8'h03;
		16'hD282: out_word = 8'hFE;
		16'hD283: out_word = 8'hE1;
		16'hD284: out_word = 8'hFD;
		16'hD285: out_word = 8'h2A;
		16'hD286: out_word = 8'h04;
		16'hD287: out_word = 8'h42;
		16'hD288: out_word = 8'hDD;
		16'hD289: out_word = 8'h7D;
		16'hD28A: out_word = 8'h17;
		16'hD28B: out_word = 8'hBD;
		16'hD28C: out_word = 8'h38;
		16'hD28D: out_word = 8'h2F;
		16'hD28E: out_word = 8'h0A;
		16'hD28F: out_word = 8'h2C;
		16'hD290: out_word = 8'h10;
		16'hD291: out_word = 8'h18;
		16'hD292: out_word = 8'hFE;
		16'hD293: out_word = 8'h02;
		16'hD294: out_word = 8'h1F;
		16'hD295: out_word = 8'h03;
		16'hD296: out_word = 8'h3D;
		16'hD297: out_word = 8'h18;
		16'hD298: out_word = 8'h17;
		16'hD299: out_word = 8'hE5;
		16'hD29A: out_word = 8'hCF;
		16'hD29B: out_word = 8'hCD;
		16'hD29C: out_word = 8'h1D;
		16'hD29D: out_word = 8'hB3;
		16'hD29E: out_word = 8'hFC;
		16'hD29F: out_word = 8'h43;
		16'hD2A0: out_word = 8'hE1;
		16'hD2A1: out_word = 8'hE8;
		16'hD2A2: out_word = 8'h38;
		16'hD2A3: out_word = 8'h41;
		16'hD2A4: out_word = 8'hE5;
		16'hD2A5: out_word = 8'hA9;
		16'hD2A6: out_word = 8'h0B;
		16'hD2A7: out_word = 8'hD3;
		16'hD2A8: out_word = 8'hE0;
		16'hD2A9: out_word = 8'h0F;
		16'hD2AA: out_word = 8'hE2;
		16'hD2AB: out_word = 8'hCD;
		16'hD2AC: out_word = 8'hD3;
		16'hD2AD: out_word = 8'hF9;
		16'hD2AE: out_word = 8'h43;
		16'hD2AF: out_word = 8'hF5;
		16'hD2B0: out_word = 8'h95;
		16'hD2B1: out_word = 8'h28;
		16'hD2B2: out_word = 8'h9E;
		16'hD2B3: out_word = 8'h2B;
		16'hD2B4: out_word = 8'hBA;
		16'hD2B5: out_word = 8'h18;
		16'hD2B6: out_word = 8'hDC;
		16'hD2B7: out_word = 8'hA7;
		16'hD2B8: out_word = 8'h52;
		16'hD2B9: out_word = 8'h79;
		16'hD2BA: out_word = 8'hF0;
		16'hD2BB: out_word = 8'hE5;
		16'hD2BC: out_word = 8'h7B;
		16'hD2BD: out_word = 8'hEF;
		16'hD2BE: out_word = 8'h3D;
		16'hD2BF: out_word = 8'h6F;
		16'hD2C0: out_word = 8'h26;
		16'hD2C1: out_word = 8'h42;
		16'hD2C2: out_word = 8'hB4;
		16'hD2C3: out_word = 8'h2F;
		16'hD2C4: out_word = 8'h81;
		16'hD2C5: out_word = 8'hE7;
		16'hD2C6: out_word = 8'h26;
		16'hD2C7: out_word = 8'hEB;
		16'hD2C8: out_word = 8'h21;
		16'hD2C9: out_word = 8'h8A;
		16'hD2CA: out_word = 8'h09;
		16'hD2CB: out_word = 8'h44;
		16'hD2CC: out_word = 8'h83;
		16'hD2CD: out_word = 8'h4D;
		16'hD2CE: out_word = 8'hD1;
		16'hD2CF: out_word = 8'hFF;
		16'hD2D0: out_word = 8'h78;
		16'hD2D1: out_word = 8'hE6;
		16'hD2D2: out_word = 8'h01;
		16'hD2D3: out_word = 8'h47;
		16'hD2D4: out_word = 8'hED;
		16'hD2D5: out_word = 8'hB0;
		16'hD2D6: out_word = 8'h21;
		16'hD2D7: out_word = 8'h58;
		16'hD2D8: out_word = 8'hE1;
		16'hD2D9: out_word = 8'h27;
		16'hD2DA: out_word = 8'hD9;
		16'hD2DB: out_word = 8'hFD;
		16'hD2DC: out_word = 8'hFA;
		16'hD2DD: out_word = 8'h3A;
		16'hD2DE: out_word = 8'h5C;
		16'hD2DF: out_word = 8'hFB;
		16'hD2E0: out_word = 8'hC3;
		16'hD2E1: out_word = 8'hFE;
		16'hD2E2: out_word = 8'h45;
		16'hD2E3: out_word = 8'hEF;
		16'hD2E4: out_word = 8'h01;
		16'hD2E5: out_word = 8'h4C;
		16'hD2E6: out_word = 8'h24;
		16'hD2E7: out_word = 8'h66;
		16'hD2E8: out_word = 8'hA7;
		16'hD2E9: out_word = 8'h3E;
		16'hD2EA: out_word = 8'h52;
		16'hD2EB: out_word = 8'h30;
		16'hD2EC: out_word = 8'h06;
		16'hD2ED: out_word = 8'h98;
		16'hD2EE: out_word = 8'h7A;
		16'hD2EF: out_word = 8'hC3;
		16'hD2F0: out_word = 8'hBE;
		16'hD2F1: out_word = 8'hA6;
		16'hD2F2: out_word = 8'hD4;
		16'hD2F3: out_word = 8'h40;
		16'hD2F4: out_word = 8'h48;
		16'hD2F5: out_word = 8'hEE;
		16'hD2F6: out_word = 8'h4E;
		16'hD2F7: out_word = 8'h92;
		16'hD2F8: out_word = 8'h4B;
		16'hD2F9: out_word = 8'hEA;
		16'hD2FA: out_word = 8'h59;
		16'hD2FB: out_word = 8'hD5;
		16'hD2FC: out_word = 8'h0A;
		16'hD2FD: out_word = 8'hF0;
		16'hD2FE: out_word = 8'h01;
		16'hD2FF: out_word = 8'h69;
		16'hD300: out_word = 8'hD7;
		16'hD301: out_word = 8'hB0;
		16'hD302: out_word = 8'hC9;
		16'hD303: out_word = 8'hCE;
		16'hD304: out_word = 8'h3A;
		16'hD305: out_word = 8'hFE;
		16'hD306: out_word = 8'h02;
		16'hD307: out_word = 8'h42;
		16'hD308: out_word = 8'hA7;
		16'hD309: out_word = 8'h20;
		16'hD30A: out_word = 8'h06;
		16'hD30B: out_word = 8'h21;
		16'hD30C: out_word = 8'hF7;
		16'hD30D: out_word = 8'hA7;
		16'hD30E: out_word = 8'h7A;
		16'hD30F: out_word = 8'hC9;
		16'hD310: out_word = 8'hB9;
		16'hD311: out_word = 8'h3D;
		16'hD312: out_word = 8'hF7;
		16'hD313: out_word = 8'hFF;
		16'hD314: out_word = 8'h40;
		16'hD315: out_word = 8'hF7;
		16'hD316: out_word = 8'h83;
		16'hD317: out_word = 8'h3B;
		16'hD318: out_word = 8'hF1;
		16'hD319: out_word = 8'h42;
		16'hD31A: out_word = 8'hC0;
		16'hD31B: out_word = 8'h41;
		16'hD31C: out_word = 8'hF4;
		16'hD31D: out_word = 8'hC6;
		16'hD31E: out_word = 8'h1E;
		16'hD31F: out_word = 8'h42;
		16'hD320: out_word = 8'h62;
		16'hD321: out_word = 8'hCE;
		16'hD322: out_word = 8'h49;
		16'hD323: out_word = 8'h21;
		16'hD324: out_word = 8'hD7;
		16'hD325: out_word = 8'h6F;
		16'hD326: out_word = 8'hC5;
		16'hD327: out_word = 8'h3F;
		16'hD328: out_word = 8'h3D;
		16'hD329: out_word = 8'hE3;
		16'hD32A: out_word = 8'h1F;
		16'hD32B: out_word = 8'hEB;
		16'hD32C: out_word = 8'h29;
		16'hD32D: out_word = 8'h29;
		16'hD32E: out_word = 8'h7F;
		16'hD32F: out_word = 8'h93;
		16'hD330: out_word = 8'hED;
		16'hD331: out_word = 8'h4A;
		16'hD332: out_word = 8'h09;
		16'hD333: out_word = 8'h7B;
		16'hD334: out_word = 8'h5A;
		16'hD335: out_word = 8'h55;
		16'hD336: out_word = 8'h4C;
		16'hD337: out_word = 8'hFE;
		16'hD338: out_word = 8'h06;
		16'hD339: out_word = 8'h00;
		16'hD33A: out_word = 8'hCD;
		16'hD33B: out_word = 8'h53;
		16'hD33C: out_word = 8'h44;
		16'hD33D: out_word = 8'h23;
		16'hD33E: out_word = 8'h4E;
		16'hD33F: out_word = 8'h37;
		16'hD340: out_word = 8'h46;
		16'hD341: out_word = 8'hED;
		16'hD342: out_word = 8'h43;
		16'hD343: out_word = 8'h49;
		16'hD344: out_word = 8'hD9;
		16'hD345: out_word = 8'h53;
		16'hD346: out_word = 8'hD9;
		16'hD347: out_word = 8'hA1;
		16'hD348: out_word = 8'hC9;
		16'hD349: out_word = 8'h5F;
		16'hD34A: out_word = 8'hE7;
		16'hD34B: out_word = 8'hF1;
		16'hD34C: out_word = 8'h51;
		16'hD34D: out_word = 8'hF5;
		16'hD34E: out_word = 8'hC5;
		16'hD34F: out_word = 8'h21;
		16'hD350: out_word = 8'hFD;
		16'hD351: out_word = 8'h42;
		16'hD352: out_word = 8'hCD;
		16'hD353: out_word = 8'h27;
		16'hD354: out_word = 8'h45;
		16'hD355: out_word = 8'h3A;
		16'hD356: out_word = 8'h4E;
		16'hD357: out_word = 8'hC1;
		16'hD358: out_word = 8'hF1;
		16'hD359: out_word = 8'h5F;
		16'hD35A: out_word = 8'h80;
		16'hD35B: out_word = 8'h00;
		16'hD35C: out_word = 8'hFF;
		16'hD35D: out_word = 8'h5E;
		16'hD35E: out_word = 8'h23;
		16'hD35F: out_word = 8'h56;
		16'hD360: out_word = 8'h18;
		16'hD361: out_word = 8'hDA;
		16'hD362: out_word = 8'hF5;
		16'hD363: out_word = 8'h62;
		16'hD364: out_word = 8'h6B;
		16'hD365: out_word = 8'h29;
		16'hD366: out_word = 8'h19;
		16'hD367: out_word = 8'h3E;
		16'hD368: out_word = 8'h96;
		16'hD369: out_word = 8'h1D;
		16'hD36A: out_word = 8'h7B;
		16'hD36B: out_word = 8'h5C;
		16'hD36C: out_word = 8'h70;
		16'hD36D: out_word = 8'hED;
		16'hD36E: out_word = 8'h42;
		16'hD36F: out_word = 8'h4A;
		16'hD370: out_word = 8'h3B;
		16'hD371: out_word = 8'h3B;
		16'hD372: out_word = 8'hF5;
		16'hD373: out_word = 8'hE5;
		16'hD374: out_word = 8'h20;
		16'hD375: out_word = 8'hD9;
		16'hD376: out_word = 8'hE7;
		16'hD377: out_word = 8'h32;
		16'hD378: out_word = 8'h09;
		16'hD379: out_word = 8'h46;
		16'hD37A: out_word = 8'h23;
		16'hD37B: out_word = 8'hF0;
		16'hD37C: out_word = 8'h7C;
		16'hD37D: out_word = 8'hFE;
		16'hD37E: out_word = 8'h42;
		16'hD37F: out_word = 8'h20;
		16'hD380: out_word = 8'h69;
		16'hD381: out_word = 8'hC5;
		16'hD382: out_word = 8'hBA;
		16'hD383: out_word = 8'h13;
		16'hD384: out_word = 8'h7B;
		16'hD385: out_word = 8'hC4;
		16'hD386: out_word = 8'h56;
		16'hD387: out_word = 8'h58;
		16'hD388: out_word = 8'h4E;
		16'hD389: out_word = 8'hF5;
		16'hD38A: out_word = 8'h1F;
		16'hD38B: out_word = 8'h30;
		16'hD38C: out_word = 8'h10;
		16'hD38D: out_word = 8'hA5;
		16'hD38E: out_word = 8'hB0;
		16'hD38F: out_word = 8'h1B;
		16'hD390: out_word = 8'h65;
		16'hD391: out_word = 8'h3F;
		16'hD392: out_word = 8'hFC;
		16'hD393: out_word = 8'h7A;
		16'hD394: out_word = 8'hE6;
		16'hD395: out_word = 8'h0F;
		16'hD396: out_word = 8'h57;
		16'hD397: out_word = 8'h18;
		16'hD398: out_word = 8'h8A;
		16'hD399: out_word = 8'h6C;
		16'hD39A: out_word = 8'h63;
		16'hD39B: out_word = 8'hFC;
		16'hD39C: out_word = 8'h78;
		16'hD39D: out_word = 8'hB1;
		16'hD39E: out_word = 8'hB2;
		16'hD39F: out_word = 8'hB3;
		16'hD3A0: out_word = 8'h20;
		16'hD3A1: out_word = 8'h13;
		16'hD3A2: out_word = 8'h93;
		16'hD3A3: out_word = 8'hF6;
		16'hD3A4: out_word = 8'hB3;
		16'hD3A5: out_word = 8'hEE;
		16'hD3A6: out_word = 8'h23;
		16'hD3A7: out_word = 8'h10;
		16'hD3A8: out_word = 8'h28;
		16'hD3A9: out_word = 8'h0B;
		16'hD3AA: out_word = 8'h34;
		16'hD3AB: out_word = 8'hE5;
		16'hD3AC: out_word = 8'hAB;
		16'hD3AD: out_word = 8'hCF;
		16'hD3AE: out_word = 8'hE1;
		16'hD3AF: out_word = 8'hC3;
		16'hD3B0: out_word = 8'hFC;
		16'hD3B1: out_word = 8'h21;
		16'hD3B2: out_word = 8'hFE;
		16'hD3B3: out_word = 8'hFF;
		16'hD3B4: out_word = 8'hC6;
		16'hD3B5: out_word = 8'hEB;
		16'hD3B6: out_word = 8'h19;
		16'hD3B7: out_word = 8'h9F;
		16'hD3B8: out_word = 8'h23;
		16'hD3B9: out_word = 8'h52;
		16'hD3BA: out_word = 8'h3A;
		16'hD3BB: out_word = 8'h04;
		16'hD3BC: out_word = 8'h42;
		16'hD3BD: out_word = 8'h18;
		16'hD3BE: out_word = 8'hBA;
		16'hD3BF: out_word = 8'h08;
		16'hD3C0: out_word = 8'h42;
		16'hD3C1: out_word = 8'hED;
		16'hD3C2: out_word = 8'h42;
		16'hD3C3: out_word = 8'h15;
		16'hD3C4: out_word = 8'hFF;
		16'hD3C5: out_word = 8'h14;
		16'hD3C6: out_word = 8'h0F;
		16'hD3C7: out_word = 8'h30;
		16'hD3C8: out_word = 8'hF5;
		16'hD3C9: out_word = 8'h44;
		16'hD3CA: out_word = 8'h4D;
		16'hD3CB: out_word = 8'h21;
		16'hD3CC: out_word = 8'h11;
		16'hD3CD: out_word = 8'h70;
		16'hD3CE: out_word = 8'h86;
		16'hD3CF: out_word = 8'h28;
		16'hD3D0: out_word = 8'h15;
		16'hD3D1: out_word = 8'h48;
		16'hD3D2: out_word = 8'hD9;
		16'hD3D3: out_word = 8'h67;
		16'hD3D4: out_word = 8'h4F;
		16'hD3D5: out_word = 8'h48;
		16'hD3D6: out_word = 8'h36;
		16'hD3D7: out_word = 8'h3E;
		16'hD3D8: out_word = 8'h02;
		16'hD3D9: out_word = 8'h48;
		16'hD3DA: out_word = 8'hDE;
		16'hD3DB: out_word = 8'h38;
		16'hD3DC: out_word = 8'hC6;
		16'hD3DD: out_word = 8'h5F;
		16'hD3DE: out_word = 8'h1A;
		16'hD3DF: out_word = 8'h53;
		16'hD3E0: out_word = 8'hA1;
		16'hD3E1: out_word = 8'hDE;
		16'hD3E2: out_word = 8'hC9;
		16'hD3E3: out_word = 8'h7E;
		16'hD3E4: out_word = 8'hE7;
		16'hD3E5: out_word = 8'h23;
		16'hD3E6: out_word = 8'h93;
		16'hD3E7: out_word = 8'h5F;
		16'hD3E8: out_word = 8'hFC;
		16'hD3E9: out_word = 8'h9A;
		16'hD3EA: out_word = 8'h57;
		16'hD3EB: out_word = 8'h38;
		16'hD3EC: out_word = 8'hFC;
		16'hD3ED: out_word = 8'h99;
		16'hD3EE: out_word = 8'h4F;
		16'hD3EF: out_word = 8'h1A;
		16'hD3F0: out_word = 8'h98;
		16'hD3F1: out_word = 8'h47;
		16'hD3F2: out_word = 8'h52;
		16'hD3F3: out_word = 8'hF0;
		16'hD3F4: out_word = 8'h83;
		16'hD3F5: out_word = 8'hF0;
		16'hD3F6: out_word = 8'h8A;
		16'hD3F7: out_word = 8'h93;
		16'hD3F8: out_word = 8'hF0;
		16'hD3F9: out_word = 8'h89;
		16'hD3FA: out_word = 8'hF0;
		16'hD3FB: out_word = 8'h88;
		16'hD3FC: out_word = 8'h38;
		16'hD3FD: out_word = 8'hF0;
		16'hD3FE: out_word = 8'hEB;
		16'hD3FF: out_word = 8'h09;
		16'hD400: out_word = 8'hC8;
		16'hD401: out_word = 8'h64;
		16'hD402: out_word = 8'h54;
		16'hD403: out_word = 8'hA5;
		16'hD404: out_word = 8'h7D;
		16'hD405: out_word = 8'h84;
		16'hD406: out_word = 8'h40;
		16'hD407: out_word = 8'hE5;
		16'hD408: out_word = 8'h3E;
		16'hD409: out_word = 8'h01;
		16'hD40A: out_word = 8'h7F;
		16'hD40B: out_word = 8'h54;
		16'hD40C: out_word = 8'hE1;
		16'hD40D: out_word = 8'hC9;
		16'hD40E: out_word = 8'h9F;
		16'hD40F: out_word = 8'hF5;
		16'hD410: out_word = 8'hF8;
		16'hD411: out_word = 8'hD3;
		16'hD412: out_word = 8'h77;
		16'hD413: out_word = 8'hF1;
		16'hD414: out_word = 8'h08;
		16'hD415: out_word = 8'h0B;
		16'hD416: out_word = 8'h52;
		16'hD417: out_word = 8'hCD;
		16'hD418: out_word = 8'hC2;
		16'hD419: out_word = 8'h89;
		16'hD41A: out_word = 8'h45;
		16'hD41B: out_word = 8'h04;
		16'hD41C: out_word = 8'h38;
		16'hD41D: out_word = 8'hE4;
		16'hD41E: out_word = 8'h71;
		16'hD41F: out_word = 8'hFE;
		16'hD420: out_word = 8'hF3;
		16'hD421: out_word = 8'h20;
		16'hD422: out_word = 8'hF9;
		16'hD423: out_word = 8'h32;
		16'hD424: out_word = 8'h57;
		16'hD425: out_word = 8'h37;
		16'hD426: out_word = 8'hD9;
		16'hD427: out_word = 8'hB2;
		16'hD428: out_word = 8'hA9;
		16'hD429: out_word = 8'hFD;
		16'hD42A: out_word = 8'h78;
		16'hD42B: out_word = 8'hFD;
		16'hD42C: out_word = 8'hC1;
		16'hD42D: out_word = 8'hFE;
		16'hD42E: out_word = 8'h08;
		16'hD42F: out_word = 8'h3D;
		16'hD430: out_word = 8'h20;
		16'hD431: out_word = 8'hE4;
		16'hD432: out_word = 8'h3E;
		16'hD433: out_word = 8'h4C;
		16'hD434: out_word = 8'hCD;
		16'hD435: out_word = 8'h3D;
		16'hD436: out_word = 8'h45;
		16'hD437: out_word = 8'h39;
		16'hD438: out_word = 8'hE0;
		16'hD439: out_word = 8'h3C;
		16'hD43A: out_word = 8'h20;
		16'hD43B: out_word = 8'hFA;
		16'hD43C: out_word = 8'hCC;
		16'hD43D: out_word = 8'h98;
		16'hD43E: out_word = 8'h03;
		16'hD43F: out_word = 8'hCC;
		16'hD440: out_word = 8'hAF;
		16'hD441: out_word = 8'hBF;
		16'hD442: out_word = 8'h57;
		16'hD443: out_word = 8'hF1;
		16'hD444: out_word = 8'hC9;
		16'hD445: out_word = 8'hE5;
		16'hD446: out_word = 8'hD5;
		16'hD447: out_word = 8'hC6;
		16'hD448: out_word = 8'hC5;
		16'hD449: out_word = 8'hF5;
		16'hD44A: out_word = 8'hD1;
		16'hD44B: out_word = 8'h3E;
		16'hD44C: out_word = 8'h7A;
		16'hD44D: out_word = 8'hD1;
		16'hD44E: out_word = 8'hA1;
		16'hD44F: out_word = 8'hE3;
		16'hD450: out_word = 8'hCB;
		16'hD451: out_word = 8'hD1;
		16'hD452: out_word = 8'h60;
		16'hD453: out_word = 8'h47;
		16'hD454: out_word = 8'hFD;
		16'hD455: out_word = 8'hCB;
		16'hD456: out_word = 8'h77;
		16'hD457: out_word = 8'hE1;
		16'hD458: out_word = 8'hD7;
		16'hD459: out_word = 8'h20;
		16'hD45A: out_word = 8'h0A;
		16'hD45B: out_word = 8'hF8;
		16'hD45C: out_word = 8'h85;
		16'hD45D: out_word = 8'hED;
		16'hD45E: out_word = 8'h6A;
		16'hD45F: out_word = 8'h65;
		16'hD460: out_word = 8'hDE;
		16'hD461: out_word = 8'h53;
		16'hD462: out_word = 8'h1E;
		16'hD463: out_word = 8'h00;
		16'hD464: out_word = 8'hF1;
		16'hD465: out_word = 8'hE4;
		16'hD466: out_word = 8'hAD;
		16'hD467: out_word = 8'h79;
		16'hD468: out_word = 8'hCC;
		16'hD469: out_word = 8'hFD;
		16'hD46A: out_word = 8'h61;
		16'hD46B: out_word = 8'hFD;
		16'hD46C: out_word = 8'h69;
		16'hD46D: out_word = 8'hCF;
		16'hD46E: out_word = 8'hFD;
		16'hD46F: out_word = 8'h51;
		16'hD470: out_word = 8'hFD;
		16'hD471: out_word = 8'h59;
		16'hD472: out_word = 8'h3E;
		16'hD473: out_word = 8'hFF;
		16'hD474: out_word = 8'h50;
		16'hD475: out_word = 8'hAB;
		16'hD476: out_word = 8'h9B;
		16'hD477: out_word = 8'hD1;
		16'hD478: out_word = 8'h7E;
		16'hD479: out_word = 8'hC5;
		16'hD47A: out_word = 8'hD4;
		16'hD47B: out_word = 8'hE6;
		16'hD47C: out_word = 8'hAF;
		16'hD47D: out_word = 8'hE3;
		16'hD47E: out_word = 8'h6C;
		16'hD47F: out_word = 8'hFD;
		16'hD480: out_word = 8'hBA;
		16'hD481: out_word = 8'h3D;
		16'hD482: out_word = 8'h1F;
		16'hD483: out_word = 8'h92;
		16'hD484: out_word = 8'hD5;
		16'hD485: out_word = 8'h11;
		16'hD486: out_word = 8'hFF;
		16'hD487: out_word = 8'h08;
		16'hD488: out_word = 8'hDB;
		16'hD489: out_word = 8'hF8;
		16'hD48A: out_word = 8'h57;
		16'hD48B: out_word = 8'hBB;
		16'hD48C: out_word = 8'h20;
		16'hD48D: out_word = 8'h03;
		16'hD48E: out_word = 8'h15;
		16'hD48F: out_word = 8'hBC;
		16'hD490: out_word = 8'hF8;
		16'hD491: out_word = 8'hD1;
		16'hD492: out_word = 8'hC9;
		16'hD493: out_word = 8'h81;
		16'hD494: out_word = 8'h5F;
		16'hD495: out_word = 8'hCD;
		16'hD496: out_word = 8'hC2;
		16'hD497: out_word = 8'h22;
		16'hD498: out_word = 8'h46;
		16'hD499: out_word = 8'h9C;
		16'hD49A: out_word = 8'hD5;
		16'hD49B: out_word = 8'hD3;
		16'hD49C: out_word = 8'hB3;
		16'hD49D: out_word = 8'h00;
		16'hD49E: out_word = 8'h2F;
		16'hD49F: out_word = 8'hD3;
		16'hD4A0: out_word = 8'hBB;
		16'hD4A1: out_word = 8'hCD;
		16'hD4A2: out_word = 8'h54;
		16'hD4A3: out_word = 8'hC0;
		16'hD4A4: out_word = 8'h46;
		16'hD4A5: out_word = 8'h11;
		16'hD4A6: out_word = 8'h85;
		16'hD4A7: out_word = 8'h02;
		16'hD4A8: out_word = 8'h4E;
		16'hD4A9: out_word = 8'h0B;
		16'hD4AA: out_word = 8'hED;
		16'hD4AB: out_word = 8'hA2;
		16'hD4AC: out_word = 8'hFA;
		16'hD4AD: out_word = 8'h1B;
		16'hD4AE: out_word = 8'h7A;
		16'hD4AF: out_word = 8'hB3;
		16'hD4B0: out_word = 8'h20;
		16'hD4B1: out_word = 8'hF6;
		16'hD4B2: out_word = 8'h50;
		16'hD4B3: out_word = 8'h5F;
		16'hD4B4: out_word = 8'hE9;
		16'hD4B5: out_word = 8'hF2;
		16'hD4B6: out_word = 8'hE4;
		16'hD4B7: out_word = 8'h81;
		16'hD4B8: out_word = 8'hFE;
		16'hD4B9: out_word = 8'h77;
		16'hD4BA: out_word = 8'h61;
		16'hD4BB: out_word = 8'hFE;
		16'hD4BC: out_word = 8'hAB;
		16'hD4BD: out_word = 8'hAF;
		16'hD4BE: out_word = 8'hC9;
		16'hD4BF: out_word = 8'hD3;
		16'hD4C0: out_word = 8'hB3;
		16'hD4C1: out_word = 8'h3E;
		16'hD4C2: out_word = 8'h1E;
		16'hD4C3: out_word = 8'hF4;
		16'hD4C4: out_word = 8'hD9;
		16'hD4C5: out_word = 8'h78;
		16'hD4C6: out_word = 8'h85;
		16'hD4C7: out_word = 8'hF6;
		16'hD4C8: out_word = 8'h48;
		16'hD4C9: out_word = 8'h0A;
		16'hD4CA: out_word = 8'h79;
		16'hD4CB: out_word = 8'hF5;
		16'hD4CC: out_word = 8'hFA;
		16'hD4CD: out_word = 8'h7A;
		16'hD4CE: out_word = 8'hEB;
		16'hD4CF: out_word = 8'hFA;
		16'hD4D0: out_word = 8'h7B;
		16'hD4D1: out_word = 8'hC4;
		16'hD4D2: out_word = 8'hFA;
		16'hD4D3: out_word = 8'hBB;
		16'hD4D4: out_word = 8'h21;
		16'hD4D5: out_word = 8'h7F;
		16'hD4D6: out_word = 8'hC9;
		16'hD4D7: out_word = 8'hDB;
		16'hD4D8: out_word = 8'hBB;
		16'hD4D9: out_word = 8'h17;
		16'hD4DA: out_word = 8'h38;
		16'hD4DB: out_word = 8'hFB;
		16'hD4DC: out_word = 8'h72;
		16'hD4DD: out_word = 8'hFA;
		16'hD4DE: out_word = 8'h30;
		16'hD4DF: out_word = 8'hE5;
		16'hD4E0: out_word = 8'hFA;
		16'hD4E1: out_word = 8'h1F;
		16'hD4E2: out_word = 8'h31;
		16'hD4E3: out_word = 8'hF4;
		16'hD4E4: out_word = 8'hC5;
		16'hD4E5: out_word = 8'hD5;
		16'hD4E6: out_word = 8'hFF;
		16'hD4E7: out_word = 8'h08;
		16'hD4E8: out_word = 8'h78;
		16'hD4E9: out_word = 8'h59;
		16'hD4EA: out_word = 8'h01;
		16'hD4EB: out_word = 8'hD0;
		16'hD4EC: out_word = 8'hFF;
		16'hD4ED: out_word = 8'hA6;
		16'hD4EE: out_word = 8'hF6;
		16'hD4EF: out_word = 8'h78;
		16'hD4F0: out_word = 8'h0E;
		16'hD4F1: out_word = 8'hB0;
		16'hD4F2: out_word = 8'h61;
		16'hD4F3: out_word = 8'h5A;
		16'hD4F4: out_word = 8'hD1;
		16'hD4F5: out_word = 8'hC8;
		16'hD4F6: out_word = 8'h90;
		16'hD4F7: out_word = 8'h52;
		16'hD4F8: out_word = 8'h92;
		16'hD4F9: out_word = 8'h70;
		16'hD4FA: out_word = 8'hF7;
		16'hD4FB: out_word = 8'h05;
		16'hD4FC: out_word = 8'h50;
		16'hD4FD: out_word = 8'h3B;
		16'hD4FE: out_word = 8'hEF;
		16'hD4FF: out_word = 8'hF0;
		16'hD500: out_word = 8'h3E;
		16'hD501: out_word = 8'h20;
		16'hD502: out_word = 8'h87;
		16'hD503: out_word = 8'hFA;
		16'hD504: out_word = 8'h98;
		16'hD505: out_word = 8'hE6;
		16'hD506: out_word = 8'h88;
		16'hD507: out_word = 8'hC8;
		16'hD508: out_word = 8'hFE;
		16'hD509: out_word = 8'h08;
		16'hD50A: out_word = 8'h68;
		16'hD50B: out_word = 8'hA7;
		16'hD50C: out_word = 8'h69;
		16'hD50D: out_word = 8'h40;
		16'hD50E: out_word = 8'h0E;
		16'hD50F: out_word = 8'hF1;
		16'hD510: out_word = 8'h10;
		16'hD511: out_word = 8'hED;
		16'hD512: out_word = 8'h58;
		16'hD513: out_word = 8'h0C;
		16'hD514: out_word = 8'h7E;
		16'hD515: out_word = 8'h50;
		16'hD516: out_word = 8'h0D;
		16'hD517: out_word = 8'h73;
		16'hD518: out_word = 8'h23;
		16'hD519: out_word = 8'h72;
		16'hD51A: out_word = 8'h33;
		16'hD51B: out_word = 8'h1C;
		16'hD51C: out_word = 8'h1B;
		16'hD51D: out_word = 8'hF6;
		16'hD51E: out_word = 8'h5C;
		16'hD51F: out_word = 8'hD5;
		16'hD520: out_word = 8'hD2;
		16'hD521: out_word = 8'hC5;
		16'hD522: out_word = 8'h80;
		16'hD523: out_word = 8'h5D;
		16'hD524: out_word = 8'h9E;
		16'hD525: out_word = 8'h50;
		16'hD526: out_word = 8'hC4;
		16'hD527: out_word = 8'hD1;
		16'hD528: out_word = 8'hC1;
		16'hD529: out_word = 8'hAF;
		16'hD52A: out_word = 8'h9F;
		16'hD52B: out_word = 8'h91;
		16'hD52C: out_word = 8'hCD;
		16'hD52D: out_word = 8'h2B;
		16'hD52E: out_word = 8'h47;
		16'hD52F: out_word = 8'h08;
		16'hD530: out_word = 8'h06;
		16'hD531: out_word = 8'h92;
		16'hD532: out_word = 8'hFF;
		16'hD533: out_word = 8'hA9;
		16'hD534: out_word = 8'h42;
		16'hD535: out_word = 8'h00;
		16'hD536: out_word = 8'hB1;
		16'hD537: out_word = 8'h56;
		16'hD538: out_word = 8'h5E;
		16'hD539: out_word = 8'hA9;
		16'hD53A: out_word = 8'h8B;
		16'hD53B: out_word = 8'hF7;
		16'hD53C: out_word = 8'hF5;
		16'hD53D: out_word = 8'hE4;
		16'hD53E: out_word = 8'h11;
		16'hD53F: out_word = 8'hD8;
		16'hD540: out_word = 8'hF8;
		16'hD541: out_word = 8'hA6;
		16'hD542: out_word = 8'h1A;
		16'hD543: out_word = 8'h42;
		16'hD544: out_word = 8'h77;
		16'hD545: out_word = 8'hEE;
		16'hD546: out_word = 8'h77;
		16'hD547: out_word = 8'h23;
		16'hD548: out_word = 8'h43;
		16'hD549: out_word = 8'h98;
		16'hD54A: out_word = 8'hFA;
		16'hD54B: out_word = 8'h44;
		16'hD54C: out_word = 8'hF4;
		16'hD54D: out_word = 8'h49;
		16'hD54E: out_word = 8'hAA;
		16'hD54F: out_word = 8'hCB;
		16'hD550: out_word = 8'hB4;
		16'hD551: out_word = 8'h44;
		16'hD552: out_word = 8'hF5;
		16'hD553: out_word = 8'h9D;
		16'hD554: out_word = 8'hCE;
		16'hD555: out_word = 8'hF9;
		16'hD556: out_word = 8'hF1;
		16'hD557: out_word = 8'hF3;
		16'hD558: out_word = 8'hB8;
		16'hD559: out_word = 8'hD1;
		16'hD55A: out_word = 8'hBF;
		16'hD55B: out_word = 8'hB9;
		16'hD55C: out_word = 8'h50;
		16'hD55D: out_word = 8'hFC;
		16'hD55E: out_word = 8'h59;
		16'hD55F: out_word = 8'h08;
		16'hD560: out_word = 8'h01;
		16'hD561: out_word = 8'hBE;
		16'hD562: out_word = 8'hFE;
		16'hD563: out_word = 8'h7A;
		16'hD564: out_word = 8'hA7;
		16'hD565: out_word = 8'h30;
		16'hD566: out_word = 8'h9E;
		16'hD567: out_word = 8'h06;
		16'hD568: out_word = 8'hFD;
		16'hD569: out_word = 8'h7B;
		16'hD56A: out_word = 8'h48;
		16'hD56B: out_word = 8'hFA;
		16'hD56C: out_word = 8'hD1;
		16'hD56D: out_word = 8'h3B;
		16'hD56E: out_word = 8'hFC;
		16'hD56F: out_word = 8'h7A;
		16'hD570: out_word = 8'h97;
		16'hD571: out_word = 8'hF3;
		16'hD572: out_word = 8'hFB;
		16'hD573: out_word = 8'h02;
		16'hD574: out_word = 8'hF3;
		16'hD575: out_word = 8'h3F;
		16'hD576: out_word = 8'h74;
		16'hD577: out_word = 8'hE5;
		16'hD578: out_word = 8'h21;
		16'hD579: out_word = 8'hF0;
		16'hD57A: out_word = 8'h3F;
		16'hD57B: out_word = 8'hE3;
		16'hD57C: out_word = 8'hE6;
		16'hD57D: out_word = 8'hC3;
		16'hD57E: out_word = 8'h2F;
		16'hD57F: out_word = 8'h3D;
		16'hD580: out_word = 8'hF8;
		16'hD581: out_word = 8'hF3;
		16'hD582: out_word = 8'hF4;
		16'hD583: out_word = 8'hF8;
		16'hD584: out_word = 8'hDD;
		16'hD585: out_word = 8'h0F;
		16'hD586: out_word = 8'h2E;
		16'hD587: out_word = 8'h68;
		16'hD588: out_word = 8'hCD;
		16'hD589: out_word = 8'hB2;
		16'hD58A: out_word = 8'h8B;
		16'hD58B: out_word = 8'h79;
		16'hD58C: out_word = 8'h8F;
		16'hD58D: out_word = 8'hF8;
		16'hD58E: out_word = 8'h62;
		16'hD58F: out_word = 8'h21;
		16'hD590: out_word = 8'h00;
		16'hD591: out_word = 8'hF8;
		16'hD592: out_word = 8'h11;
		16'hD593: out_word = 8'hB8;
		16'hD594: out_word = 8'hC0;
		16'hD595: out_word = 8'h01;
		16'hD596: out_word = 8'h55;
		16'hD597: out_word = 8'h08;
		16'hD598: out_word = 8'hDF;
		16'hD599: out_word = 8'h4B;
		16'hD59A: out_word = 8'h72;
		16'hD59B: out_word = 8'h67;
		16'hD59C: out_word = 8'h11;
		16'hD59D: out_word = 8'h3A;
		16'hD59E: out_word = 8'hF4;
		16'hD59F: out_word = 8'h5C;
		16'hD5A0: out_word = 8'h01;
		16'hD5A1: out_word = 8'hBC;
		16'hD5A2: out_word = 8'h00;
		16'hD5A3: out_word = 8'hF5;
		16'hD5A4: out_word = 8'hE1;
		16'hD5A5: out_word = 8'h76;
		16'hD5A6: out_word = 8'h75;
		16'hD5A7: out_word = 8'hE5;
		16'hD5A8: out_word = 8'h70;
		16'hD5A9: out_word = 8'h73;
		16'hD5AA: out_word = 8'h3D;
		16'hD5AB: out_word = 8'h5C;
		16'hD5AC: out_word = 8'h3F;
		16'hD5AD: out_word = 8'h58;
		16'hD5AE: out_word = 8'hFF;
		16'hD5AF: out_word = 8'hF9;
		16'hD5B0: out_word = 8'h11;
		16'hD5B1: out_word = 8'h08;
		16'hD5B2: out_word = 8'h3E;
		16'hD5B3: out_word = 8'hF4;
		16'hD5B4: out_word = 8'h01;
		16'hD5B5: out_word = 8'hA8;
		16'hD5B6: out_word = 8'h00;
		16'hD5B7: out_word = 8'hEB;
		16'hD5B8: out_word = 8'hEB;
		16'hD5B9: out_word = 8'h0E;
		16'hD5BA: out_word = 8'h3E;
		16'hD5BB: out_word = 8'h71;
		16'hD5BC: out_word = 8'hC0;
		16'hD5BD: out_word = 8'h03;
		16'hD5BE: out_word = 8'h13;
		16'hD5BF: out_word = 8'h0C;
		16'hD5C0: out_word = 8'hE3;
		16'hD5C1: out_word = 8'h1B;
		16'hD5C2: out_word = 8'h03;
		16'hD5C3: out_word = 8'hBF;
		16'hD5C4: out_word = 8'hD1;
		16'hD5C5: out_word = 8'hF0;
		16'hD5C6: out_word = 8'h5C;
		16'hD5C7: out_word = 8'hC3;
		16'hD5C8: out_word = 8'h3E;
		16'hD5C9: out_word = 8'h07;
		16'hD5CA: out_word = 8'hB2;
		16'hD5CB: out_word = 8'h60;
		16'hD5CC: out_word = 8'h6F;
		16'hD5CD: out_word = 8'hC2;
		16'hD5CE: out_word = 8'h63;
		16'hD5CF: out_word = 8'hCD;
		16'hD5D0: out_word = 8'h70;
		16'hD5D1: out_word = 8'h21;
		16'hD5D2: out_word = 8'hE2;
		16'hD5D3: out_word = 8'hBA;
		16'hD5D4: out_word = 8'h97;
		16'hD5D5: out_word = 8'h11;
		16'hD5D6: out_word = 8'hB4;
		16'hD5D7: out_word = 8'hA2;
		16'hD5D8: out_word = 8'hB7;
		16'hD5D9: out_word = 8'hAF;
		16'hD5DA: out_word = 8'hCE;
		16'hD5DB: out_word = 8'h43;
		16'hD5DC: out_word = 8'hC5;
		16'hD5DD: out_word = 8'hD3;
		16'hD5DE: out_word = 8'hFE;
		16'hD5DF: out_word = 8'h27;
		16'hD5E0: out_word = 8'h32;
		16'hD5E1: out_word = 8'h8A;
		16'hD5E2: out_word = 8'h6C;
		16'hD5E3: out_word = 8'hE5;
		16'hD5E4: out_word = 8'hCD;
		16'hD5E5: out_word = 8'h46;
		16'hD5E6: out_word = 8'h63;
		16'hD5E7: out_word = 8'hC2;
		16'hD5E8: out_word = 8'h39;
		16'hD5E9: out_word = 8'hF8;
		16'hD5EA: out_word = 8'hC3;
		16'hD5EB: out_word = 8'h62;
		16'hD5EC: out_word = 8'h60;
		16'hD5ED: out_word = 8'h7D;
		16'hD5EE: out_word = 8'hE6;
		16'hD5EF: out_word = 8'h07;
		16'hD5F0: out_word = 8'h18;
		16'hD5F1: out_word = 8'h0D;
		16'hD5F2: out_word = 8'hFB;
		16'hD5F3: out_word = 8'h09;
		16'hD5F4: out_word = 8'h1C;
		16'hD5F5: out_word = 8'h08;
		16'hD5F6: out_word = 8'hC3;
		16'hD5F7: out_word = 8'hFB;
		16'hD5F8: out_word = 8'h0B;
		16'hD5F9: out_word = 8'h9F;
		16'hD5FA: out_word = 8'h03;
		16'hD5FB: out_word = 8'hFB;
		16'hD5FC: out_word = 8'h0D;
		16'hD5FD: out_word = 8'h22;
		16'hD5FE: out_word = 8'hF6;
		16'hD5FF: out_word = 8'h6B;
		16'hD600: out_word = 8'hF1;
		16'hD601: out_word = 8'hF3;
		16'hD602: out_word = 8'h3E;
		16'hD603: out_word = 8'hF7;
		16'hD604: out_word = 8'hCD;
		16'hD605: out_word = 8'h69;
		16'hD606: out_word = 8'h63;
		16'hD607: out_word = 8'hC4;
		16'hD608: out_word = 8'h54;
		16'hD609: out_word = 8'hFD;
		16'hD60A: out_word = 8'h5D;
		16'hD60B: out_word = 8'h13;
		16'hD60C: out_word = 8'h01;
		16'hD60D: out_word = 8'hFF;
		16'hD60E: out_word = 8'h0F;
		16'hD60F: out_word = 8'h75;
		16'hD610: out_word = 8'h3F;
		16'hD611: out_word = 8'hB8;
		16'hD612: out_word = 8'hF2;
		16'hD613: out_word = 8'h6B;
		16'hD614: out_word = 8'h11;
		16'hD615: out_word = 8'hE1;
		16'hD616: out_word = 8'hC8;
		16'hD617: out_word = 8'h0E;
		16'hD618: out_word = 8'h94;
		16'hD619: out_word = 8'h1C;
		16'hD61A: out_word = 8'hF6;
		16'hD61B: out_word = 8'hCC;
		16'hD61C: out_word = 8'hF4;
		16'hD61D: out_word = 8'h3E;
		16'hD61E: out_word = 8'h80;
		16'hD61F: out_word = 8'hD3;
		16'hD620: out_word = 8'h33;
		16'hD621: out_word = 8'hF9;
		16'hD622: out_word = 8'h9A;
		16'hD623: out_word = 8'hDD;
		16'hD624: out_word = 8'h8D;
		16'hD625: out_word = 8'h69;
		16'hD626: out_word = 8'h73;
		16'hD627: out_word = 8'h51;
		16'hD628: out_word = 8'hC3;
		16'hD629: out_word = 8'hF7;
		16'hD62A: out_word = 8'h75;
		16'hD62B: out_word = 8'hF6;
		16'hD62C: out_word = 8'h6A;
		16'hD62D: out_word = 8'h73;
		16'hD62E: out_word = 8'h47;
		16'hD62F: out_word = 8'h18;
		16'hD630: out_word = 8'h07;
		16'hD631: out_word = 8'h33;
		16'hD632: out_word = 8'hF7;
		16'hD633: out_word = 8'h25;
		16'hD634: out_word = 8'hA3;
		16'hD635: out_word = 8'h98;
		16'hD636: out_word = 8'hF8;
		16'hD637: out_word = 8'h7E;
		16'hD638: out_word = 8'hED;
		16'hD639: out_word = 8'h7B;
		16'hD63A: out_word = 8'h64;
		16'hD63B: out_word = 8'h60;
		16'hD63C: out_word = 8'h3C;
		16'hD63D: out_word = 8'h3C;
		16'hD63E: out_word = 8'h63;
		16'hD63F: out_word = 8'hFB;
		16'hD640: out_word = 8'h41;
		16'hD641: out_word = 8'hA0;
		16'hD642: out_word = 8'h85;
		16'hD643: out_word = 8'hFB;
		16'hD644: out_word = 8'h30;
		16'hD645: out_word = 8'h62;
		16'hD646: out_word = 8'h3E;
		16'hD647: out_word = 8'hFF;
		16'hD648: out_word = 8'h31;
		16'hD649: out_word = 8'h8D;
		16'hD64A: out_word = 8'hCD;
		16'hD64B: out_word = 8'hD3;
		16'hD64C: out_word = 8'h03;
		16'hD64D: out_word = 8'h63;
		16'hD64E: out_word = 8'h1D;
		16'hD64F: out_word = 8'hF3;
		16'hD650: out_word = 8'hAF;
		16'hD651: out_word = 8'h4B;
		16'hD652: out_word = 8'h9D;
		16'hD653: out_word = 8'hC7;
		16'hD654: out_word = 8'h43;
		16'hD655: out_word = 8'hF4;
		16'hD656: out_word = 8'h51;
		16'hD657: out_word = 8'hF9;
		16'hD658: out_word = 8'hC2;
		16'hD659: out_word = 8'h52;
		16'hD65A: out_word = 8'h7E;
		16'hD65B: out_word = 8'hCE;
		16'hD65C: out_word = 8'h26;
		16'hD65D: out_word = 8'h86;
		16'hD65E: out_word = 8'hF9;
		16'hD65F: out_word = 8'h9F;
		16'hD660: out_word = 8'h65;
		16'hD661: out_word = 8'hE4;
		16'hD662: out_word = 8'hA8;
		16'hD663: out_word = 8'h83;
		16'hD664: out_word = 8'hC0;
		16'hD665: out_word = 8'h97;
		16'hD666: out_word = 8'hD7;
		16'hD667: out_word = 8'hCE;
		16'hD668: out_word = 8'h50;
		16'hD669: out_word = 8'h76;
		16'hD66A: out_word = 8'h74;
		16'hD66B: out_word = 8'h18;
		16'hD66C: out_word = 8'h02;
		16'hD66D: out_word = 8'h25;
		16'hD66E: out_word = 8'h17;
		16'hD66F: out_word = 8'h12;
		16'hD670: out_word = 8'hF7;
		16'hD671: out_word = 8'hC5;
		16'hD672: out_word = 8'hF3;
		16'hD673: out_word = 8'h47;
		16'hD674: out_word = 8'h33;
		16'hD675: out_word = 8'h4F;
		16'hD676: out_word = 8'hDB;
		16'hD677: out_word = 8'h39;
		16'hD678: out_word = 8'hFE;
		16'hD679: out_word = 8'h15;
		16'hD67A: out_word = 8'h28;
		16'hD67B: out_word = 8'h89;
		16'hD67C: out_word = 8'h34;
		16'hD67D: out_word = 8'h12;
		16'hD67E: out_word = 8'h12;
		16'hD67F: out_word = 8'h30;
		16'hD680: out_word = 8'h04;
		16'hD681: out_word = 8'h10;
		16'hD682: out_word = 8'h0A;
		16'hD683: out_word = 8'h2C;
		16'hD684: out_word = 8'hD7;
		16'hD685: out_word = 8'h22;
		16'hD686: out_word = 8'hED;
		16'hD687: out_word = 8'h79;
		16'hD688: out_word = 8'h31;
		16'hD689: out_word = 8'h3B;
		16'hD68A: out_word = 8'hEB;
		16'hD68B: out_word = 8'h42;
		16'hD68C: out_word = 8'hD5;
		16'hD68D: out_word = 8'h1D;
		16'hD68E: out_word = 8'h7F;
		16'hD68F: out_word = 8'hFF;
		16'hD690: out_word = 8'h10;
		16'hD691: out_word = 8'hDE;
		16'hD692: out_word = 8'hF9;
		16'hD693: out_word = 8'h4F;
		16'hD694: out_word = 8'hE6;
		16'hD695: out_word = 8'hC7;
		16'hD696: out_word = 8'hC8;
		16'hD697: out_word = 8'h17;
		16'hD698: out_word = 8'h07;
		16'hD699: out_word = 8'h79;
		16'hD69A: out_word = 8'hFE;
		16'hD69B: out_word = 8'h20;
		16'hD69C: out_word = 8'h02;
		16'hD69D: out_word = 8'hD6;
		16'hD69E: out_word = 8'h38;
		16'hD69F: out_word = 8'h3D;
		16'hD6A0: out_word = 8'h18;
		16'hD6A1: out_word = 8'hBA;
		16'hD6A2: out_word = 8'h7E;
		16'hD6A3: out_word = 8'hB6;
		16'hD6A4: out_word = 8'hD0;
		16'hD6A5: out_word = 8'hE5;
		16'hD6A6: out_word = 8'hCD;
		16'hD6A7: out_word = 8'h12;
		16'hD6A8: out_word = 8'h8E;
		16'hD6A9: out_word = 8'h17;
		16'hD6AA: out_word = 8'h7C;
		16'hD6AB: out_word = 8'hE1;
		16'hD6AC: out_word = 8'hA7;
		16'hD6AD: out_word = 8'hFF;
		16'hD6AE: out_word = 8'h20;
		16'hD6AF: out_word = 8'h0B;
		16'hD6B0: out_word = 8'hE5;
		16'hD6B1: out_word = 8'hEB;
		16'hD6B2: out_word = 8'h21;
		16'hD6B3: out_word = 8'hC0;
		16'hD6B4: out_word = 8'h76;
		16'hD6B5: out_word = 8'h01;
		16'hD6B6: out_word = 8'hD7;
		16'hD6B7: out_word = 8'h50;
		16'hD6B8: out_word = 8'h00;
		16'hD6B9: out_word = 8'h0D;
		16'hD6BA: out_word = 8'h13;
		16'hD6BB: out_word = 8'h7F;
		16'hD6BC: out_word = 8'h41;
		16'hD6BD: out_word = 8'hA9;
		16'hD6BE: out_word = 8'h27;
		16'hD6BF: out_word = 8'hDB;
		16'hD6C0: out_word = 8'h08;
		16'hD6C1: out_word = 8'hC3;
		16'hD6C2: out_word = 8'h11;
		16'hD6C3: out_word = 8'h02;
		16'hD6C4: out_word = 8'h5E;
		16'hD6C5: out_word = 8'h69;
		16'hD6C6: out_word = 8'hDF;
		16'hD6C7: out_word = 8'h3E;
		16'hD6C8: out_word = 8'hE0;
		16'hD6C9: out_word = 8'hEB;
		16'hD6CA: out_word = 8'h69;
		16'hD6CB: out_word = 8'h51;
		16'hD6CC: out_word = 8'h23;
		16'hD6CD: out_word = 8'hD9;
		16'hD6CE: out_word = 8'h6A;
		16'hD6CF: out_word = 8'h3E;
		16'hD6D0: out_word = 8'h30;
		16'hD6D1: out_word = 8'hEE;
		16'hD6D2: out_word = 8'hB1;
		16'hD6D3: out_word = 8'h08;
		16'hD6D4: out_word = 8'h0F;
		16'hD6D5: out_word = 8'h57;
		16'hD6D6: out_word = 8'h67;
		16'hD6D7: out_word = 8'hAF;
		16'hD6D8: out_word = 8'h99;
		16'hD6D9: out_word = 8'h68;
		16'hD6DA: out_word = 8'h3E;
		16'hD6DB: out_word = 8'h86;
		16'hD6DC: out_word = 8'hB2;
		16'hD6DD: out_word = 8'hF3;
		16'hD6DE: out_word = 8'h7D;
		16'hD6DF: out_word = 8'h86;
		16'hD6E0: out_word = 8'hE3;
		16'hD6E1: out_word = 8'hFE;
		16'hD6E2: out_word = 8'hC9;
		16'hD6E3: out_word = 8'h3A;
		16'hD6E4: out_word = 8'h50;
		16'hD6E5: out_word = 8'h6C;
		16'hD6E6: out_word = 8'h32;
		16'hD6E7: out_word = 8'h30;
		16'hD6E8: out_word = 8'h77;
		16'hD6E9: out_word = 8'h6E;
		16'hD6EA: out_word = 8'hA0;
		16'hD6EB: out_word = 8'h0E;
		16'hD6EC: out_word = 8'hFA;
		16'hD6ED: out_word = 8'hDA;
		16'hD6EE: out_word = 8'hFF;
		16'hD6EF: out_word = 8'hE5;
		16'hD6F0: out_word = 8'h3A;
		16'hD6F1: out_word = 8'h08;
		16'hD6F2: out_word = 8'h5C;
		16'hD6F3: out_word = 8'hFF;
		16'hD6F4: out_word = 8'hD6;
		16'hD6F5: out_word = 8'h31;
		16'hD6F6: out_word = 8'hFE;
		16'hD6F7: out_word = 8'h04;
		16'hD6F8: out_word = 8'h30;
		16'hD6F9: out_word = 8'h27;
		16'hD6FA: out_word = 8'h32;
		16'hD6FB: out_word = 8'h3D;
		16'hD6FC: out_word = 8'hA5;
		16'hD6FD: out_word = 8'h77;
		16'hD6FE: out_word = 8'h25;
		16'hD6FF: out_word = 8'h3E;
		16'hD700: out_word = 8'h6C;
		16'hD701: out_word = 8'hDC;
		16'hD702: out_word = 8'h0F;
		16'hD703: out_word = 8'h01;
		16'hD704: out_word = 8'h05;
		16'hD705: out_word = 8'h40;
		16'hD706: out_word = 8'hD5;
		16'hD707: out_word = 8'h07;
		16'hD708: out_word = 8'h13;
		16'hD709: out_word = 8'h3D;
		16'hD70A: out_word = 8'hB4;
		16'hD70B: out_word = 8'hD1;
		16'hD70C: out_word = 8'h68;
		16'hD70D: out_word = 8'hF3;
		16'hD70E: out_word = 8'h06;
		16'hD70F: out_word = 8'h40;
		16'hD710: out_word = 8'hF4;
		16'hD711: out_word = 8'hED;
		16'hD712: out_word = 8'h7D;
		16'hD713: out_word = 8'h7A;
		16'hD714: out_word = 8'h7A;
		16'hD715: out_word = 8'hFE;
		16'hD716: out_word = 8'hA0;
		16'hD717: out_word = 8'h20;
		16'hD718: out_word = 8'hDF;
		16'hD719: out_word = 8'hDF;
		16'hD71A: out_word = 8'hC2;
		16'hD71B: out_word = 8'hC5;
		16'hD71C: out_word = 8'h8A;
		16'hD71D: out_word = 8'h85;
		16'hD71E: out_word = 8'hBB;
		16'hD71F: out_word = 8'h0E;
		16'hD720: out_word = 8'hF5;
		16'hD721: out_word = 8'h64;
		16'hD722: out_word = 8'hC9;
		16'hD723: out_word = 8'hF0;
		16'hD724: out_word = 8'h9E;
		16'hD725: out_word = 8'h69;
		16'hD726: out_word = 8'hA1;
		16'hD727: out_word = 8'hC9;
		16'hD728: out_word = 8'hE8;
		16'hD729: out_word = 8'hD3;
		16'hD72A: out_word = 8'h06;
		16'hD72B: out_word = 8'h08;
		16'hD72C: out_word = 8'h4B;
		16'hD72D: out_word = 8'hF3;
		16'hD72E: out_word = 8'hCD;
		16'hD72F: out_word = 8'hFE;
		16'hD730: out_word = 8'h5D;
		16'hD731: out_word = 8'h77;
		16'hD732: out_word = 8'h3E;
		16'hD733: out_word = 8'hA0;
		16'hD734: out_word = 8'h32;
		16'hD735: out_word = 8'h6F;
		16'hD736: out_word = 8'hE8;
		16'hD737: out_word = 8'h04;
		16'hD738: out_word = 8'h6E;
		16'hD739: out_word = 8'h50;
		16'hD73A: out_word = 8'h3F;
		16'hD73B: out_word = 8'h0C;
		16'hD73C: out_word = 8'h01;
		16'hD73D: out_word = 8'hC8;
		16'hD73E: out_word = 8'h00;
		16'hD73F: out_word = 8'hC5;
		16'hD740: out_word = 8'hCD;
		16'hD741: out_word = 8'hD6;
		16'hD742: out_word = 8'h73;
		16'hD743: out_word = 8'hE8;
		16'hD744: out_word = 8'h3D;
		16'hD745: out_word = 8'hFA;
		16'hD746: out_word = 8'hFE;
		16'hD747: out_word = 8'h3E;
		16'hD748: out_word = 8'h08;
		16'hD749: out_word = 8'hC1;
		16'hD74A: out_word = 8'h05;
		16'hD74B: out_word = 8'hF6;
		16'hD74C: out_word = 8'h99;
		16'hD74D: out_word = 8'h5E;
		16'hD74E: out_word = 8'hEA;
		16'hD74F: out_word = 8'h10;
		16'hD750: out_word = 8'hAF;
		16'hD751: out_word = 8'h03;
		16'hD752: out_word = 8'hDB;
		16'hD753: out_word = 8'hF0;
		16'hD754: out_word = 8'hCF;
		16'hD755: out_word = 8'hCB;
		16'hD756: out_word = 8'h7F;
		16'hD757: out_word = 8'h73;
		16'hD758: out_word = 8'hE6;
		16'hD759: out_word = 8'hE9;
		16'hD75A: out_word = 8'hFE;
		16'hD75B: out_word = 8'h85;
		16'hD75C: out_word = 8'h40;
		16'hD75D: out_word = 8'hD1;
		16'hD75E: out_word = 8'hDC;
		16'hD75F: out_word = 8'hC3;
		16'hD760: out_word = 8'h00;
		16'hD761: out_word = 8'hE9;
		16'hD762: out_word = 8'h20;
		16'hD763: out_word = 8'h23;
		16'hD764: out_word = 8'h94;
		16'hD765: out_word = 8'hC8;
		16'hD766: out_word = 8'hDE;
		16'hD767: out_word = 8'h02;
		16'hD768: out_word = 8'hB0;
		16'hD769: out_word = 8'h05;
		16'hD76A: out_word = 8'hAF;
		16'hD76B: out_word = 8'hC8;
		16'hD76C: out_word = 8'hF9;
		16'hD76D: out_word = 8'h90;
		16'hD76E: out_word = 8'h2E;
		16'hD76F: out_word = 8'h4D;
		16'hD770: out_word = 8'hFA;
		16'hD771: out_word = 8'h70;
		16'hD772: out_word = 8'hEB;
		16'hD773: out_word = 8'h03;
		16'hD774: out_word = 8'h17;
		16'hD775: out_word = 8'hF8;
		16'hD776: out_word = 8'hCA;
		16'hD777: out_word = 8'hEF;
		16'hD778: out_word = 8'h18;
		16'hD779: out_word = 8'h14;
		16'hD77A: out_word = 8'hF8;
		16'hD77B: out_word = 8'h1A;
		16'hD77C: out_word = 8'hC4;
		16'hD77D: out_word = 8'h77;
		16'hD77E: out_word = 8'hF3;
		16'hD77F: out_word = 8'hF2;
		16'hD780: out_word = 8'h06;
		16'hD781: out_word = 8'h30;
		16'hD782: out_word = 8'hA8;
		16'hD783: out_word = 8'h4B;
		16'hD784: out_word = 8'h40;
		16'hD785: out_word = 8'hA8;
		16'hD786: out_word = 8'hB1;
		16'hD787: out_word = 8'h01;
		16'hD788: out_word = 8'h10;
		16'hD789: out_word = 8'h30;
		16'hD78A: out_word = 8'hED;
		16'hD78B: out_word = 8'hA2;
		16'hD78C: out_word = 8'hE9;
		16'hD78D: out_word = 8'h11;
		16'hD78E: out_word = 8'hFB;
		16'hD78F: out_word = 8'hC1;
		16'hD790: out_word = 8'hCC;
		16'hD791: out_word = 8'h10;
		16'hD792: out_word = 8'hF2;
		16'hD793: out_word = 8'hFD;
		16'hD794: out_word = 8'hE9;
		16'hD795: out_word = 8'hFF;
		16'hD796: out_word = 8'h71;
		16'hD797: out_word = 8'h65;
		16'hD798: out_word = 8'hE8;
		16'hD799: out_word = 8'hCB;
		16'hD79A: out_word = 8'h5F;
		16'hD79B: out_word = 8'hC0;
		16'hD79C: out_word = 8'h18;
		16'hD79D: out_word = 8'hF8;
		16'hD79E: out_word = 8'hA7;
		16'hD79F: out_word = 8'hF5;
		16'hD7A0: out_word = 8'h7F;
		16'hD7A1: out_word = 8'hF1;
		16'hD7A2: out_word = 8'h01;
		16'hD7A3: out_word = 8'hF0;
		16'hD7A4: out_word = 8'h71;
		16'hD7A5: out_word = 8'hBA;
		16'hD7A6: out_word = 8'h3D;
		16'hD7A7: out_word = 8'hED;
		16'hD7A8: out_word = 8'h07;
		16'hD7A9: out_word = 8'hD0;
		16'hD7AA: out_word = 8'h18;
		16'hD7AB: out_word = 8'hF9;
		16'hD7AC: out_word = 8'h0A;
		16'hD7AD: out_word = 8'hEF;
		16'hD7AE: out_word = 8'hF0;
		16'hD7AF: out_word = 8'hE7;
		16'hD7B0: out_word = 8'h31;
		16'hD7B1: out_word = 8'hC9;
		16'hD7B2: out_word = 8'h3E;
		16'hD7B3: out_word = 8'hB0;
		16'hD7B4: out_word = 8'h2B;
		16'hD7B5: out_word = 8'h93;
		16'hD7B6: out_word = 8'hA0;
		16'hD7B7: out_word = 8'h21;
		16'hD7B8: out_word = 8'h21;
		16'hD7B9: out_word = 8'h8A;
		16'hD7BA: out_word = 8'h6A;
		16'hD7BB: out_word = 8'h40;
		16'hD7BC: out_word = 8'hAF;
		16'hD7BD: out_word = 8'hE9;
		16'hD7BE: out_word = 8'hEC;
		16'hD7BF: out_word = 8'hFB;
		16'hD7C0: out_word = 8'h06;
		16'hD7C1: out_word = 8'hF0;
		16'hD7C2: out_word = 8'h1E;
		16'hD7C3: out_word = 8'h76;
		16'hD7C4: out_word = 8'h10;
		16'hD7C5: out_word = 8'hFD;
		16'hD7C6: out_word = 8'h3F;
		16'hD7C7: out_word = 8'h3D;
		16'hD7C8: out_word = 8'hE9;
		16'hD7C9: out_word = 8'h01;
		16'hD7CA: out_word = 8'h14;
		16'hD7CB: out_word = 8'hEB;
		16'hD7CC: out_word = 8'hB7;
		16'hD7CD: out_word = 8'hF3;
		16'hD7CE: out_word = 8'hED;
		16'hD7CF: out_word = 8'h42;
		16'hD7D0: out_word = 8'hC2;
		16'hD7D1: out_word = 8'h76;
		16'hD7D2: out_word = 8'h99;
		16'hD7D3: out_word = 8'hD7;
		16'hD7D4: out_word = 8'hE2;
		16'hD7D5: out_word = 8'hE9;
		16'hD7D6: out_word = 8'hCD;
		16'hD7D7: out_word = 8'h70;
		16'hD7D8: out_word = 8'h85;
		16'hD7D9: out_word = 8'hE3;
		16'hD7DA: out_word = 8'h71;
		16'hD7DB: out_word = 8'hFA;
		16'hD7DC: out_word = 8'hE3;
		16'hD7DD: out_word = 8'hE3;
		16'hD7DE: out_word = 8'h25;
		16'hD7DF: out_word = 8'h9D;
		16'hD7E0: out_word = 8'h37;
		16'hD7E1: out_word = 8'hF1;
		16'hD7E2: out_word = 8'hFB;
		16'hD7E3: out_word = 8'h11;
		16'hD7E4: out_word = 8'hF1;
		16'hD7E5: out_word = 8'hC7;
		16'hD7E6: out_word = 8'h11;
		16'hD7E7: out_word = 8'h82;
		16'hD7E8: out_word = 8'hD3;
		16'hD7E9: out_word = 8'h6C;
		16'hD7EA: out_word = 8'h6B;
		16'hD7EB: out_word = 8'h81;
		16'hD7EC: out_word = 8'h73;
		16'hD7ED: out_word = 8'h4C;
		16'hD7EE: out_word = 8'h43;
		16'hD7EF: out_word = 8'hEF;
		16'hD7F0: out_word = 8'hD1;
		16'hD7F1: out_word = 8'h01;
		16'hD7F2: out_word = 8'hFF;
		16'hD7F3: out_word = 8'h60;
		16'hD7F4: out_word = 8'h7E;
		16'hD7F5: out_word = 8'hC6;
		16'hD7F6: out_word = 8'hF6;
		16'hD7F7: out_word = 8'h6F;
		16'hD7F8: out_word = 8'h16;
		16'hD7F9: out_word = 8'h87;
		16'hD7FA: out_word = 8'hCD;
		16'hD7FB: out_word = 8'h9E;
		16'hD7FC: out_word = 8'h0E;
		16'hD7FD: out_word = 8'hBC;
		16'hD7FE: out_word = 8'hA2;
		16'hD7FF: out_word = 8'h80;
		16'hD800: out_word = 8'h09;
		16'hD801: out_word = 8'h91;
		16'hD802: out_word = 8'hF9;
		16'hD803: out_word = 8'hE5;
		16'hD804: out_word = 8'h60;
		16'hD805: out_word = 8'h21;
		16'hD806: out_word = 8'hC0;
		16'hD807: out_word = 8'h11;
		16'hD808: out_word = 8'h04;
		16'hD809: out_word = 8'h2F;
		16'hD80A: out_word = 8'h0A;
		16'hD80B: out_word = 8'h1A;
		16'hD80C: out_word = 8'hED;
		16'hD80D: out_word = 8'hA1;
		16'hD80E: out_word = 8'hFF;
		16'hD80F: out_word = 8'h20;
		16'hD810: out_word = 8'h18;
		16'hD811: out_word = 8'h13;
		16'hD812: out_word = 8'hEA;
		16'hD813: out_word = 8'hDF;
		16'hD814: out_word = 8'hE8;
		16'hD815: out_word = 8'hE1;
		16'hD816: out_word = 8'h0E;
		16'hD817: out_word = 8'hBC;
		16'hD818: out_word = 8'h06;
		16'hD819: out_word = 8'hE7;
		16'hD81A: out_word = 8'h56;
		16'hD81B: out_word = 8'h7E;
		16'hD81C: out_word = 8'hF0;
		16'hD81D: out_word = 8'h77;
		16'hD81E: out_word = 8'h11;
		16'hD81F: out_word = 8'hFB;
		16'hD820: out_word = 8'hF0;
		16'hD821: out_word = 8'h21;
		16'hD822: out_word = 8'h04;
		16'hD823: out_word = 8'h75;
		16'hD824: out_word = 8'hC9;
		16'hD825: out_word = 8'hE1;
		16'hD826: out_word = 8'hAF;
		16'hD827: out_word = 8'h73;
		16'hD828: out_word = 8'h2B;
		16'hD829: out_word = 8'h78;
		16'hD82A: out_word = 8'hB1;
		16'hD82B: out_word = 8'h20;
		16'hD82C: out_word = 8'hFF;
		16'hD82D: out_word = 8'h02;
		16'hD82E: out_word = 8'h24;
		16'hD82F: out_word = 8'h6F;
		16'hD830: out_word = 8'h09;
		16'hD831: out_word = 8'h7C;
		16'hD832: out_word = 8'hFE;
		16'hD833: out_word = 8'h40;
		16'hD834: out_word = 8'h30;
		16'hD835: out_word = 8'hF9;
		16'hD836: out_word = 8'hC9;
		16'hD837: out_word = 8'hC7;
		16'hD838: out_word = 8'hD5;
		16'hD839: out_word = 8'h11;
		16'hD83A: out_word = 8'hF1;
		16'hD83B: out_word = 8'hBD;
		16'hD83C: out_word = 8'hAF;
		16'hD83D: out_word = 8'h04;
		16'hD83E: out_word = 8'h75;
		16'hD83F: out_word = 8'hFD;
		16'hD840: out_word = 8'hD1;
		16'hD841: out_word = 8'h38;
		16'hD842: out_word = 8'h03;
		16'hD843: out_word = 8'hAC;
		16'hD844: out_word = 8'h7A;
		16'hD845: out_word = 8'hEB;
		16'hD846: out_word = 8'h37;
		16'hD847: out_word = 8'hEB;
		16'hD848: out_word = 8'h21;
		16'hD849: out_word = 8'h08;
		16'hD84A: out_word = 8'h04;
		16'hD84B: out_word = 8'h37;
		16'hD84C: out_word = 8'hDE;
		16'hD84D: out_word = 8'hFB;
		16'hD84E: out_word = 8'h0C;
		16'hD84F: out_word = 8'h06;
		16'hD850: out_word = 8'h08;
		16'hD851: out_word = 8'hA0;
		16'hD852: out_word = 8'hE2;
		16'hD853: out_word = 8'hC0;
		16'hD854: out_word = 8'h21;
		16'hD855: out_word = 8'hF4;
		16'hD856: out_word = 8'h7C;
		16'hD857: out_word = 8'h34;
		16'hD858: out_word = 8'h2B;
		16'hD859: out_word = 8'h28;
		16'hD85A: out_word = 8'hFC;
		16'hD85B: out_word = 8'hE1;
		16'hD85C: out_word = 8'hC4;
		16'hD85D: out_word = 8'h0F;
		16'hD85E: out_word = 8'hF0;
		16'hD85F: out_word = 8'hBB;
		16'hD860: out_word = 8'hC9;
		16'hD861: out_word = 8'hFD;
		16'hD862: out_word = 8'hD5;
		16'hD863: out_word = 8'h6B;
		16'hD864: out_word = 8'hE8;
		16'hD865: out_word = 8'h6F;
		16'hD866: out_word = 8'h7D;
		16'hD867: out_word = 8'hC7;
		16'hD868: out_word = 8'h3B;
		16'hD869: out_word = 8'hF9;
		16'hD86A: out_word = 8'h67;
		16'hD86B: out_word = 8'hC9;
		16'hD86C: out_word = 8'hC5;
		16'hD86D: out_word = 8'h46;
		16'hD86E: out_word = 8'h62;
		16'hD86F: out_word = 8'hC1;
		16'hD870: out_word = 8'h03;
		16'hD871: out_word = 8'hED;
		16'hD872: out_word = 8'h2F;
		16'hD873: out_word = 8'hE5;
		16'hD874: out_word = 8'hB9;
		16'hD875: out_word = 8'hE0;
		16'hD876: out_word = 8'hEA;
		16'hD877: out_word = 8'h77;
		16'hD878: out_word = 8'h81;
		16'hD879: out_word = 8'h23;
		16'hD87A: out_word = 8'h11;
		16'hD87B: out_word = 8'h7A;
		16'hD87C: out_word = 8'hF8;
		16'hD87D: out_word = 8'hC1;
		16'hD87E: out_word = 8'h7A;
		16'hD87F: out_word = 8'h76;
		16'hD880: out_word = 8'hEA;
		16'hD881: out_word = 8'h59;
		16'hD882: out_word = 8'hE9;
		16'hD883: out_word = 8'h3F;
		16'hD884: out_word = 8'hCD;
		16'hD885: out_word = 8'hE8;
		16'hD886: out_word = 8'h9B;
		16'hD887: out_word = 8'hCD;
		16'hD888: out_word = 8'hBE;
		16'hD889: out_word = 8'hFF;
		16'hD88A: out_word = 8'hBF;
		16'hD88B: out_word = 8'hA9;
		16'hD88C: out_word = 8'hA0;
		16'hD88D: out_word = 8'h77;
		16'hD88E: out_word = 8'hC7;
		16'hD88F: out_word = 8'hFF;
		16'hD890: out_word = 8'hE8;
		16'hD891: out_word = 8'hC5;
		16'hD892: out_word = 8'h23;
		16'hD893: out_word = 8'h7E;
		16'hD894: out_word = 8'hD9;
		16'hD895: out_word = 8'h90;
		16'hD896: out_word = 8'hF0;
		16'hD897: out_word = 8'h2B;
		16'hD898: out_word = 8'h11;
		16'hD899: out_word = 8'hC9;
		16'hD89A: out_word = 8'h23;
		16'hD89B: out_word = 8'hF8;
		16'hD89C: out_word = 8'h23;
		16'hD89D: out_word = 8'h9D;
		16'hD89E: out_word = 8'h9F;
		16'hD89F: out_word = 8'hEA;
		16'hD8A0: out_word = 8'hC9;
		16'hD8A1: out_word = 8'hC1;
		16'hD8A2: out_word = 8'h8A;
		16'hD8A3: out_word = 8'h2E;
		16'hD8A4: out_word = 8'hEF;
		16'hD8A5: out_word = 8'h51;
		16'hD8A6: out_word = 8'h08;
		16'hD8A7: out_word = 8'hE1;
		16'hD8A8: out_word = 8'hA5;
		16'hD8A9: out_word = 8'h79;
		16'hD8AA: out_word = 8'hE0;
		16'hD8AB: out_word = 8'hFF;
		16'hD8AC: out_word = 8'h9D;
		16'hD8AD: out_word = 8'hE1;
		16'hD8AE: out_word = 8'h20;
		16'hD8AF: out_word = 8'h0F;
		16'hD8B0: out_word = 8'h13;
		16'hD8B1: out_word = 8'hF3;
		16'hD8B2: out_word = 8'h52;
		16'hD8B3: out_word = 8'h28;
		16'hD8B4: out_word = 8'hF4;
		16'hD8B5: out_word = 8'hE6;
		16'hD8B6: out_word = 8'hD7;
		16'hD8B7: out_word = 8'h7B;
		16'hD8B8: out_word = 8'hE6;
		16'hD8B9: out_word = 8'h18;
		16'hD8BA: out_word = 8'hDC;
		16'hD8BB: out_word = 8'h5D;
		16'hD8BC: out_word = 8'h22;
		16'hD8BD: out_word = 8'h5F;
		16'hD8BE: out_word = 8'hF6;
		16'hD8BF: out_word = 8'h9F;
		16'hD8C0: out_word = 8'hC3;
		16'hD8C1: out_word = 8'hDE;
		16'hD8C2: out_word = 8'h41;
		16'hD8C3: out_word = 8'h55;
		16'hD8C4: out_word = 8'h54;
		16'hD8C5: out_word = 8'h4F;
		16'hD8C6: out_word = 8'h89;
		16'hD8C7: out_word = 8'h52;
		16'hD8C8: out_word = 8'h4E;
		16'hD8C9: out_word = 8'hEC;
		16'hD8CA: out_word = 8'h2E;
		16'hD8CB: out_word = 8'h5A;
		16'hD8CC: out_word = 8'h58;
		16'hD8CD: out_word = 8'hAB;
		16'hD8CE: out_word = 8'hCD;
		16'hD8CF: out_word = 8'h8E;
		16'hD8D0: out_word = 8'hBB;
		16'hD8D1: out_word = 8'hFD;
		16'hD8D2: out_word = 8'hB0;
		16'hD8D3: out_word = 8'hB2;
		16'hD8D4: out_word = 8'hF4;
		16'hD8D5: out_word = 8'h28;
		16'hD8D6: out_word = 8'hDA;
		16'hD8D7: out_word = 8'hC9;
		16'hD8D8: out_word = 8'hEE;
		16'hD8D9: out_word = 8'hFC;
		16'hD8DA: out_word = 8'h43;
		16'hD8DB: out_word = 8'h78;
		16'hD8DC: out_word = 8'hF6;
		16'hD8DD: out_word = 8'hA2;
		16'hD8DE: out_word = 8'hC4;
		16'hD8DF: out_word = 8'hFC;
		16'hD8E0: out_word = 8'h6B;
		16'hD8E1: out_word = 8'h6C;
		16'hD8E2: out_word = 8'hA1;
		16'hD8E3: out_word = 8'h7A;
		16'hD8E4: out_word = 8'hDF;
		16'hD8E5: out_word = 8'hC0;
		16'hD8E6: out_word = 8'hC3;
		16'hD8E7: out_word = 8'h76;
		16'hD8E8: out_word = 8'hE8;
		16'hD8E9: out_word = 8'hDD;
		16'hD8EA: out_word = 8'hCB;
		16'hD8EB: out_word = 8'h87;
		16'hD8EC: out_word = 8'h08;
		16'hD8ED: out_word = 8'h21;
		16'hD8EE: out_word = 8'hFD;
		16'hD8EF: out_word = 8'h01;
		16'hD8F0: out_word = 8'h80;
		16'hD8F1: out_word = 8'h06;
		16'hD8F2: out_word = 8'hFF;
		16'hD8F3: out_word = 8'h28;
		16'hD8F4: out_word = 8'h04;
		16'hD8F5: out_word = 8'h77;
		16'hD8F6: out_word = 8'h97;
		16'hD8F7: out_word = 8'h45;
		16'hD8F8: out_word = 8'h7C;
		16'hD8F9: out_word = 8'hF1;
		16'hD8FA: out_word = 8'h32;
		16'hD8FB: out_word = 8'h53;
		16'hD8FC: out_word = 8'h7B;
		16'hD8FD: out_word = 8'h7D;
		16'hD8FE: out_word = 8'h22;
		16'hD8FF: out_word = 8'h60;
		16'hD900: out_word = 8'h40;
		16'hD901: out_word = 8'h78;
		16'hD902: out_word = 8'h80;
		16'hD903: out_word = 8'h87;
		16'hD904: out_word = 8'h0C;
		16'hD905: out_word = 8'h6F;
		16'hD906: out_word = 8'h1E;
		16'hD907: out_word = 8'hDD;
		16'hD908: out_word = 8'h6E;
		16'hD909: out_word = 8'h00;
		16'hD90A: out_word = 8'h2E;
		16'hD90B: out_word = 8'h66;
		16'hD90C: out_word = 8'h01;
		16'hD90D: out_word = 8'h16;
		16'hD90E: out_word = 8'h4E;
		16'hD90F: out_word = 8'h02;
		16'hD910: out_word = 8'h16;
		16'hD911: out_word = 8'h46;
		16'hD912: out_word = 8'h03;
		16'hD913: out_word = 8'h17;
		16'hD914: out_word = 8'h7E;
		16'hD915: out_word = 8'h04;
		16'hD916: out_word = 8'hCD;
		16'hD917: out_word = 8'hD3;
		16'hD918: out_word = 8'h1E;
		16'hD919: out_word = 8'h7B;
		16'hD91A: out_word = 8'hD0;
		16'hD91B: out_word = 8'h6E;
		16'hD91C: out_word = 8'h28;
		16'hD91D: out_word = 8'h8F;
		16'hD91E: out_word = 8'h21;
		16'hD91F: out_word = 8'h5F;
		16'hD920: out_word = 8'hC7;
		16'hD921: out_word = 8'h7C;
		16'hD922: out_word = 8'h35;
		16'hD923: out_word = 8'hCF;
		16'hD924: out_word = 8'hDD;
		16'hD925: out_word = 8'hE5;
		16'hD926: out_word = 8'hE7;
		16'hD927: out_word = 8'h00;
		16'hD928: out_word = 8'h06;
		16'hD929: out_word = 8'h08;
		16'hD92A: out_word = 8'h38;
		16'hD92B: out_word = 8'hDC;
		16'hD92C: out_word = 8'h01;
		16'hD92D: out_word = 8'h26;
		16'hD92E: out_word = 8'h2B;
		16'hD92F: out_word = 8'hBA;
		16'hD930: out_word = 8'h35;
		16'hD931: out_word = 8'hF6;
		16'hD932: out_word = 8'h29;
		16'hD933: out_word = 8'h7C;
		16'hD934: out_word = 8'hFF;
		16'hD935: out_word = 8'hEB;
		16'hD936: out_word = 8'hDD;
		16'hD937: out_word = 8'h19;
		16'hD938: out_word = 8'hCD;
		16'hD939: out_word = 8'h05;
		16'hD93A: out_word = 8'hD2;
		16'hD93B: out_word = 8'hDB;
		16'hD93C: out_word = 8'hE1;
		16'hD93D: out_word = 8'hD9;
		16'hD93E: out_word = 8'h7E;
		16'hD93F: out_word = 8'h5B;
		16'hD940: out_word = 8'hD9;
		16'hD941: out_word = 8'h08;
		16'hD942: out_word = 8'hDE;
		16'hD943: out_word = 8'h1A;
		16'hD944: out_word = 8'h1B;
		16'hD945: out_word = 8'h86;
		16'hD946: out_word = 8'h02;
		16'hD947: out_word = 8'hB0;
		16'hD948: out_word = 8'h54;
		16'hD949: out_word = 8'hE3;
		16'hD94A: out_word = 8'hDD;
		16'hD94B: out_word = 8'h8D;
		16'hD94C: out_word = 8'hD5;
		16'hD94D: out_word = 8'hDC;
		16'hD94E: out_word = 8'hD9;
		16'hD94F: out_word = 8'h7E;
		16'hD950: out_word = 8'h00;
		16'hD951: out_word = 8'h87;
		16'hD952: out_word = 8'hF9;
		16'hD953: out_word = 8'hFF;
		16'hD954: out_word = 8'h3C;
		16'hD955: out_word = 8'h57;
		16'hD956: out_word = 8'h32;
		16'hD957: out_word = 8'hA2;
		16'hD958: out_word = 8'h8B;
		16'hD959: out_word = 8'h8A;
		16'hD95A: out_word = 8'h84;
		16'hD95B: out_word = 8'h89;
		16'hD95C: out_word = 8'hD8;
		16'hD95D: out_word = 8'hF2;
		16'hD95E: out_word = 8'h5F;
		16'hD95F: out_word = 8'hF2;
		16'hD960: out_word = 8'hED;
		16'hD961: out_word = 8'h53;
		16'hD962: out_word = 8'h03;
		16'hD963: out_word = 8'h7E;
		16'hD964: out_word = 8'hF5;
		16'hD965: out_word = 8'h22;
		16'hD966: out_word = 8'h40;
		16'hD967: out_word = 8'hF5;
		16'hD968: out_word = 8'h32;
		16'hD969: out_word = 8'hB9;
		16'hD96A: out_word = 8'h7D;
		16'hD96B: out_word = 8'h90;
		16'hD96C: out_word = 8'hC4;
		16'hD96D: out_word = 8'hD1;
		16'hD96E: out_word = 8'hE2;
		16'hD96F: out_word = 8'h7C;
		16'hD970: out_word = 8'h64;
		16'hD971: out_word = 8'h39;
		16'hD972: out_word = 8'hF6;
		16'hD973: out_word = 8'h66;
		16'hD974: out_word = 8'h20;
		16'hD975: out_word = 8'h09;
		16'hD976: out_word = 8'h92;
		16'hD977: out_word = 8'h9F;
		16'hD978: out_word = 8'h0D;
		16'hD979: out_word = 8'h6E;
		16'hD97A: out_word = 8'h0E;
		16'hD97B: out_word = 8'hCD;
		16'hD97C: out_word = 8'h5C;
		16'hD97D: out_word = 8'h7D;
		16'hD97E: out_word = 8'hFF;
		16'hD97F: out_word = 8'h22;
		16'hD980: out_word = 8'h6C;
		16'hD981: out_word = 8'h61;
		16'hD982: out_word = 8'hC9;
		16'hD983: out_word = 8'h06;
		16'hD984: out_word = 8'h18;
		16'hD985: out_word = 8'h11;
		16'hD986: out_word = 8'h00;
		16'hD987: out_word = 8'hA6;
		16'hD988: out_word = 8'h40;
		16'hD989: out_word = 8'hB1;
		16'hD98A: out_word = 8'h0E;
		16'hD98B: out_word = 8'h08;
		16'hD98C: out_word = 8'hEE;
		16'hD98D: out_word = 8'hFC;
		16'hD98E: out_word = 8'h83;
		16'hD98F: out_word = 8'h14;
		16'hD990: out_word = 8'h0D;
		16'hD991: out_word = 8'h20;
		16'hD992: out_word = 8'hF8;
		16'hD993: out_word = 8'h3E;
		16'hD994: out_word = 8'h5F;
		16'hD995: out_word = 8'h83;
		16'hD996: out_word = 8'h5F;
		16'hD997: out_word = 8'h38;
		16'hD998: out_word = 8'h04;
		16'hD999: out_word = 8'hF5;
		16'hD99A: out_word = 8'h7A;
		16'hD99B: out_word = 8'hD6;
		16'hD99C: out_word = 8'h08;
		16'hD99D: out_word = 8'h57;
		16'hD99E: out_word = 8'hF3;
		16'hD99F: out_word = 8'hB0;
		16'hD9A0: out_word = 8'hD4;
		16'hD9A1: out_word = 8'h06;
		16'hD9A2: out_word = 8'h3F;
		16'hD9A3: out_word = 8'hD4;
		16'hD9A4: out_word = 8'h07;
		16'hD9A5: out_word = 8'h87;
		16'hD9A6: out_word = 8'h16;
		16'hD9A7: out_word = 8'h00;
		16'hD9A8: out_word = 8'h5F;
		16'hD9A9: out_word = 8'hBB;
		16'hD9AA: out_word = 8'h19;
		16'hD9AB: out_word = 8'hFE;
		16'hD9AC: out_word = 8'h22;
		16'hD9AD: out_word = 8'h7D;
		16'hD9AE: out_word = 8'hB4;
		16'hD9AF: out_word = 8'hC8;
		16'hD9B0: out_word = 8'hE9;
		16'hD9B1: out_word = 8'h9F;
		16'hD9B2: out_word = 8'hB8;
		16'hD9B3: out_word = 8'h54;
		16'hD9B4: out_word = 8'h5D;
		16'hD9B5: out_word = 8'h39;
		16'hD9B6: out_word = 8'h06;
		16'hD9B7: out_word = 8'h60;
		16'hD9B8: out_word = 8'h81;
		16'hD9B9: out_word = 8'h31;
		16'hD9BA: out_word = 8'h58;
		16'hD9BB: out_word = 8'h61;
		16'hD9BC: out_word = 8'h0F;
		16'hD9BD: out_word = 8'h13;
		16'hD9BE: out_word = 8'hC1;
		16'hD9BF: out_word = 8'hD2;
		16'hD9C0: out_word = 8'h57;
		16'hD9C1: out_word = 8'h5F;
		16'hD9C2: out_word = 8'h9E;
		16'hD9C3: out_word = 8'h39;
		16'hD9C4: out_word = 8'hD4;
		16'hD9C5: out_word = 8'h5B;
		16'hD9C6: out_word = 8'h06;
		16'hD9C7: out_word = 8'h0C;
		16'hD9C8: out_word = 8'hC2;
		16'hD9C9: out_word = 8'h14;
		16'hD9CA: out_word = 8'hD2;
		16'hD9CB: out_word = 8'h0F;
		16'hD9CC: out_word = 8'hFD;
		16'hD9CD: out_word = 8'hFF;
		16'hD9CE: out_word = 8'hE6;
		16'hD9CF: out_word = 8'h07;
		16'hD9D0: out_word = 8'hD3;
		16'hD9D1: out_word = 8'hFE;
		16'hD9D2: out_word = 8'hC9;
		16'hD9D3: out_word = 8'h05;
		16'hD9D4: out_word = 8'h2B;
		16'hD9D5: out_word = 8'hE5;
		16'hD9D6: out_word = 8'h23;
		16'hD9D7: out_word = 8'h81;
		16'hD9D8: out_word = 8'h6F;
		16'hD9D9: out_word = 8'h85;
		16'hD9DA: out_word = 8'h0F;
		16'hD9DB: out_word = 8'hF9;
		16'hD9DC: out_word = 8'h93;
		16'hD9DD: out_word = 8'h1C;
		16'hD9DE: out_word = 8'h36;
		16'hD9DF: out_word = 8'hFF;
		16'hD9E0: out_word = 8'h5E;
		16'hD9E1: out_word = 8'hD7;
		16'hD9E2: out_word = 8'hFF;
		16'hD9E3: out_word = 8'h7C;
		16'hD9E4: out_word = 8'hC1;
		16'hD9E5: out_word = 8'h10;
		16'hD9E6: out_word = 8'hE8;
		16'hD9E7: out_word = 8'hC9;
		16'hD9E8: out_word = 8'hE5;
		16'hD9E9: out_word = 8'hC5;
		16'hD9EA: out_word = 8'hDD;
		16'hD9EB: out_word = 8'h17;
		16'hD9EC: out_word = 8'hF5;
		16'hD9ED: out_word = 8'h3E;
		16'hD9EE: out_word = 8'hCF;
		16'hD9EF: out_word = 8'h22;
		16'hD9F0: out_word = 8'h90;
		16'hD9F1: out_word = 8'h28;
		16'hD9F2: out_word = 8'h5F;
		16'hD9F3: out_word = 8'h7C;
		16'hD9F4: out_word = 8'hC5;
		16'hD9F5: out_word = 8'hCC;
		16'hD9F6: out_word = 8'h79;
		16'hD9F7: out_word = 8'h07;
		16'hD9F8: out_word = 8'hFF;
		16'hD9F9: out_word = 8'h3D;
		16'hD9FA: out_word = 8'h7B;
		16'hD9FB: out_word = 8'h47;
		16'hD9FC: out_word = 8'hFF;
		16'hD9FD: out_word = 8'hF2;
		16'hD9FE: out_word = 8'h6A;
		16'hD9FF: out_word = 8'h86;
		16'hDA00: out_word = 8'h26;
		16'hDA01: out_word = 8'hD7;
		16'hDA02: out_word = 8'hE6;
		16'hDA03: out_word = 8'hC3;
		16'hDA04: out_word = 8'hDF;
		16'hDA05: out_word = 8'h4D;
		16'hDA06: out_word = 8'h52;
		16'hDA07: out_word = 8'hCB;
		16'hDA08: out_word = 8'hFE;
		16'hDA09: out_word = 8'h5E;
		16'hDA0A: out_word = 8'h79;
		16'hDA0B: out_word = 8'hC4;
		16'hDA0C: out_word = 8'h56;
		16'hDA0D: out_word = 8'h01;
		16'hDA0E: out_word = 8'h79;
		16'hDA0F: out_word = 8'h34;
		16'hDA10: out_word = 8'hF1;
		16'hDA11: out_word = 8'hEB;
		16'hDA12: out_word = 8'h36;
		16'hDA13: out_word = 8'h80;
		16'hDA14: out_word = 8'h23;
		16'hDA15: out_word = 8'h68;
		16'hDA16: out_word = 8'h00;
		16'hDA17: out_word = 8'hBA;
		16'hDA18: out_word = 8'hF7;
		16'hDA19: out_word = 8'hBC;
		16'hDA1A: out_word = 8'h36;
		16'hDA1B: out_word = 8'h01;
		16'hDA1C: out_word = 8'h10;
		16'hDA1D: out_word = 8'hB4;
		16'hDA1E: out_word = 8'hE1;
		16'hDA1F: out_word = 8'h5E;
		16'hDA20: out_word = 8'hE5;
		16'hDA21: out_word = 8'h14;
		16'hDA22: out_word = 8'hE4;
		16'hDA23: out_word = 8'hB5;
		16'hDA24: out_word = 8'hFF;
		16'hDA25: out_word = 8'h7B;
		16'hDA26: out_word = 8'hE7;
		16'hDA27: out_word = 8'hED;
		16'hDA28: out_word = 8'hA0;
		16'hDA29: out_word = 8'hC1;
		16'hDA2A: out_word = 8'hDD;
		16'hDA2B: out_word = 8'h53;
		16'hDA2C: out_word = 8'hE7;
		16'hDA2D: out_word = 8'h3C;
		16'hDA2E: out_word = 8'hE8;
		16'hDA2F: out_word = 8'h75;
		16'hDA30: out_word = 8'h73;
		16'hDA31: out_word = 8'h81;
		16'hDA32: out_word = 8'h5F;
		16'hDA33: out_word = 8'hF9;
		16'hDA34: out_word = 8'hA7;
		16'hDA35: out_word = 8'h1F;
		16'hDA36: out_word = 8'hFF;
		16'hDA37: out_word = 8'hFF;
		16'hDA38: out_word = 8'hE6;
		16'hDA39: out_word = 8'h0F;
		16'hDA3A: out_word = 8'hF6;
		16'hDA3B: out_word = 8'h50;
		16'hDA3C: out_word = 8'h57;
		16'hDA3D: out_word = 8'hEB;
		16'hDA3E: out_word = 8'hD1;
		16'hDA3F: out_word = 8'h43;
		16'hDA40: out_word = 8'hD2;
		16'hDA41: out_word = 8'hF1;
		16'hDA42: out_word = 8'hE5;
		16'hDA43: out_word = 8'hE1;
		16'hDA44: out_word = 8'h77;
		16'hDA45: out_word = 8'hD5;
		16'hDA46: out_word = 8'hE0;
		16'hDA47: out_word = 8'hE1;
		16'hDA48: out_word = 8'hFC;
		16'hDA49: out_word = 8'h11;
		16'hDA4A: out_word = 8'h20;
		16'hDA4B: out_word = 8'h00;
		16'hDA4C: out_word = 8'h19;
		16'hDA4D: out_word = 8'h10;
		16'hDA4E: out_word = 8'hED;
		16'hDA4F: out_word = 8'h9A;
		16'hDA50: out_word = 8'hC1;
		16'hDA51: out_word = 8'hF6;
		16'hDA52: out_word = 8'hC9;
		16'hDA53: out_word = 8'h2F;
		16'hDA54: out_word = 8'h61;
		16'hDA55: out_word = 8'hF9;
		16'hDA56: out_word = 8'h33;
		16'hDA57: out_word = 8'h2C;
		16'hDA58: out_word = 8'hCD;
		16'hDA59: out_word = 8'hA1;
		16'hDA5A: out_word = 8'h7C;
		16'hDA5B: out_word = 8'hCF;
		16'hDA5C: out_word = 8'hB9;
		16'hDA5D: out_word = 8'h10;
		16'hDA5E: out_word = 8'h3F;
		16'hDA5F: out_word = 8'h11;
		16'hDA60: out_word = 8'h79;
		16'hDA61: out_word = 8'hC2;
		16'hDA62: out_word = 8'h3E;
		16'hDA63: out_word = 8'hAA;
		16'hDA64: out_word = 8'hCD;
		16'hDA65: out_word = 8'h13;
		16'hDA66: out_word = 8'h7C;
		16'hDA67: out_word = 8'h11;
		16'hDA68: out_word = 8'h10;
		16'hDA69: out_word = 8'h4D;
		16'hDA6A: out_word = 8'hA1;
		16'hDA6B: out_word = 8'hD7;
		16'hDA6C: out_word = 8'hE6;
		16'hDA6D: out_word = 8'h1E;
		16'hDA6E: out_word = 8'hD7;
		16'hDA6F: out_word = 8'hD8;
		16'hDA70: out_word = 8'hC3;
		16'hDA71: out_word = 8'h7E;
		16'hDA72: out_word = 8'h02;
		16'hDA73: out_word = 8'hFB;
		16'hDA74: out_word = 8'h86;
		16'hDA75: out_word = 8'h01;
		16'hDA76: out_word = 8'hD6;
		16'hDA77: out_word = 8'h03;
		16'hDA78: out_word = 8'h6F;
		16'hDA79: out_word = 8'hD7;
		16'hDA7A: out_word = 8'hD3;
		16'hDA7B: out_word = 8'h00;
		16'hDA7C: out_word = 8'h28;
		16'hDA7D: out_word = 8'hD3;
		16'hDA7E: out_word = 8'h01;
		16'hDA7F: out_word = 8'hCB;
		16'hDA80: out_word = 8'hE5;
		16'hDA81: out_word = 8'hD3;
		16'hDA82: out_word = 8'h11;
		16'hDA83: out_word = 8'hCD;
		16'hDA84: out_word = 8'hD3;
		16'hDA85: out_word = 8'hF0;
		16'hDA86: out_word = 8'hFF;
		16'hDA87: out_word = 8'hBB;
		16'hDA88: out_word = 8'hD3;
		16'hDA89: out_word = 8'hE5;
		16'hDA8A: out_word = 8'hD5;
		16'hDA8B: out_word = 8'h4F;
		16'hDA8C: out_word = 8'h96;
		16'hDA8D: out_word = 8'hD1;
		16'hDA8E: out_word = 8'hE1;
		16'hDA8F: out_word = 8'h24;
		16'hDA90: out_word = 8'h14;
		16'hDA91: out_word = 8'h61;
		16'hDA92: out_word = 8'hE8;
		16'hDA93: out_word = 8'hF7;
		16'hDA94: out_word = 8'hE5;
		16'hDA95: out_word = 8'hB5;
		16'hDA96: out_word = 8'h18;
		16'hDA97: out_word = 8'hFE;
		16'hDA98: out_word = 8'h4F;
		16'hDA99: out_word = 8'h87;
		16'hDA9A: out_word = 8'h8F;
		16'hDA9B: out_word = 8'hFE;
		16'hDA9C: out_word = 8'hC9;
		16'hDA9D: out_word = 8'h3E;
		16'hDA9E: out_word = 8'h20;
		16'hDA9F: out_word = 8'hDD;
		16'hDAA0: out_word = 8'hDD;
		16'hDAA1: out_word = 8'h96;
		16'hDAA2: out_word = 8'h03;
		16'hDAA3: out_word = 8'hF5;
		16'hDAA4: out_word = 8'h80;
		16'hDAA5: out_word = 8'hE1;
		16'hDAA6: out_word = 8'h67;
		16'hDAA7: out_word = 8'h79;
		16'hDAA8: out_word = 8'h46;
		16'hDAA9: out_word = 8'h02;
		16'hDAAA: out_word = 8'h05;
		16'hDAAB: out_word = 8'hFF;
		16'hDAAC: out_word = 8'h5F;
		16'hDAAD: out_word = 8'h85;
		16'hDAAE: out_word = 8'h6F;
		16'hDAAF: out_word = 8'hE3;
		16'hDAB0: out_word = 8'h6C;
		16'hDAB1: out_word = 8'hFE;
		16'hDAB2: out_word = 8'hC9;
		16'hDAB3: out_word = 8'hFF;
		16'hDAB4: out_word = 8'h32;
		16'hDAB5: out_word = 8'hE0;
		16'hDAB6: out_word = 8'h7C;
		16'hDAB7: out_word = 8'h7D;
		16'hDAB8: out_word = 8'hE6;
		16'hDAB9: out_word = 8'h18;
		16'hDABA: out_word = 8'hF6;
		16'hDABB: out_word = 8'h40;
		16'hDABC: out_word = 8'h9A;
		16'hDABD: out_word = 8'h08;
		16'hDABE: out_word = 8'hFA;
		16'hDABF: out_word = 8'h07;
		16'hDAC0: out_word = 8'hFF;
		16'hDAC1: out_word = 8'h2F;
		16'hDAC2: out_word = 8'h84;
		16'hDAC3: out_word = 8'h6F;
		16'hDAC4: out_word = 8'h08;
		16'hDAC5: out_word = 8'hEE;
		16'hDAC6: out_word = 8'h67;
		16'hDAC7: out_word = 8'h5D;
		16'hDAC8: out_word = 8'h7C;
		16'hDAC9: out_word = 8'hFF;
		16'hDACA: out_word = 8'h26;
		16'hDACB: out_word = 8'h03;
		16'hDACC: out_word = 8'hF6;
		16'hDACD: out_word = 8'h58;
		16'hDACE: out_word = 8'hEF;
		16'hDACF: out_word = 8'h57;
		16'hDAD0: out_word = 8'h3E;
		16'hDAD1: out_word = 8'h00;
		16'hDAD2: out_word = 8'hFF;
		16'hDAD3: out_word = 8'h23;
		16'hDAD4: out_word = 8'h86;
		16'hDAD5: out_word = 8'h03;
		16'hDAD6: out_word = 8'h67;
		16'hDAD7: out_word = 8'h5F;
		16'hDAD8: out_word = 8'hD8;
		16'hDAD9: out_word = 8'hF5;
		16'hDADA: out_word = 8'hCD;
		16'hDADB: out_word = 8'hC2;
		16'hDADC: out_word = 8'h7C;
		16'hDADD: out_word = 8'hEB;
		16'hDADE: out_word = 8'hDE;
		16'hDADF: out_word = 8'hEC;
		16'hDAE0: out_word = 8'hE6;
		16'hDAE1: out_word = 8'h47;
		16'hDAE2: out_word = 8'h4F;
		16'hDAE3: out_word = 8'h2C;
		16'hDAE4: out_word = 8'h40;
		16'hDAE5: out_word = 8'h4F;
		16'hDAE6: out_word = 8'h2D;
		16'hDAE7: out_word = 8'h79;
		16'hDAE8: out_word = 8'hC6;
		16'hDAE9: out_word = 8'h28;
		16'hDAEA: out_word = 8'h87;
		16'hDAEB: out_word = 8'h77;
		16'hDAEC: out_word = 8'h3E;
		16'hDAED: out_word = 8'hD2;
		16'hDAEE: out_word = 8'h25;
		16'hDAEF: out_word = 8'hB0;
		16'hDAF0: out_word = 8'hFB;
		16'hDAF1: out_word = 8'h34;
		16'hDAF2: out_word = 8'hE5;
		16'hDAF3: out_word = 8'hFB;
		16'hDAF4: out_word = 8'h16;
		16'hDAF5: out_word = 8'h25;
		16'hDAF6: out_word = 8'hFB;
		16'hDAF7: out_word = 8'h79;
		16'hDAF8: out_word = 8'hBD;
		16'hDAF9: out_word = 8'h3F;
		16'hDAFA: out_word = 8'hFF;
		16'hDAFB: out_word = 8'hB0;
		16'hDAFC: out_word = 8'hC6;
		16'hDAFD: out_word = 8'h02;
		16'hDAFE: out_word = 8'h77;
		16'hDAFF: out_word = 8'hEB;
		16'hDB00: out_word = 8'h2D;
		16'hDB01: out_word = 8'hFC;
		16'hDB02: out_word = 8'h06;
		16'hDB03: out_word = 8'h08;
		16'hDB04: out_word = 8'hAF;
		16'hDB05: out_word = 8'h4D;
		16'hDB06: out_word = 8'h37;
		16'hDB07: out_word = 8'h17;
		16'hDB08: out_word = 8'hB5;
		16'hDB09: out_word = 8'hEC;
		16'hDB0A: out_word = 8'h7C;
		16'hDB0B: out_word = 8'hFE;
		16'hDB0C: out_word = 8'h69;
		16'hDB0D: out_word = 8'h24;
		16'hDB0E: out_word = 8'h10;
		16'hDB0F: out_word = 8'hF1;
		16'hDB10: out_word = 8'hC9;
		16'hDB11: out_word = 8'h49;
		16'hDB12: out_word = 8'h7C;
		16'hDB13: out_word = 8'hDF;
		16'hDB14: out_word = 8'hFF;
		16'hDB15: out_word = 8'hC0;
		16'hDB16: out_word = 8'h7D;
		16'hDB17: out_word = 8'hC6;
		16'hDB18: out_word = 8'h20;
		16'hDB19: out_word = 8'h6F;
		16'hDB1A: out_word = 8'hD8;
		16'hDB1B: out_word = 8'h7C;
		16'hDB1C: out_word = 8'hD6;
		16'hDB1D: out_word = 8'h3A;
		16'hDB1E: out_word = 8'h99;
		16'hDB1F: out_word = 8'hC9;
		16'hDB20: out_word = 8'h25;
		16'hDB21: out_word = 8'h52;
		16'hDB22: out_word = 8'hF1;
		16'hDB23: out_word = 8'hFE;
		16'hDB24: out_word = 8'hEF;
		16'hDB25: out_word = 8'hD6;
		16'hDB26: out_word = 8'hE4;
		16'hDB27: out_word = 8'hEF;
		16'hDB28: out_word = 8'hC6;
		16'hDB29: out_word = 8'hA7;
		16'hDB2A: out_word = 8'hEF;
		16'hDB2B: out_word = 8'h53;
		16'hDB2C: out_word = 8'h85;
		16'hDB2D: out_word = 8'h6F;
		16'hDB2E: out_word = 8'hD0;
		16'hDB2F: out_word = 8'hD1;
		16'hDB30: out_word = 8'h18;
		16'hDB31: out_word = 8'hF4;
		16'hDB32: out_word = 8'hEF;
		16'hDB33: out_word = 8'h3F;
		16'hDB34: out_word = 8'hF9;
		16'hDB35: out_word = 8'hDC;
		16'hDB36: out_word = 8'h7E;
		16'hDB37: out_word = 8'h23;
		16'hDB38: out_word = 8'hA7;
		16'hDB39: out_word = 8'hC8;
		16'hDB3A: out_word = 8'hCD;
		16'hDB3B: out_word = 8'hFF;
		16'hDB3C: out_word = 8'h65;
		16'hDB3D: out_word = 8'h7D;
		16'hDB3E: out_word = 8'h18;
		16'hDB3F: out_word = 8'hF7;
		16'hDB40: out_word = 8'hFE;
		16'hDB41: out_word = 8'h20;
		16'hDB42: out_word = 8'hD2;
		16'hDB43: out_word = 8'hF5;
		16'hDB44: out_word = 8'h04;
		16'hDB45: out_word = 8'h38;
		16'hDB46: out_word = 8'h03;
		16'hDB47: out_word = 8'h5F;
		16'hDB48: out_word = 8'h1C;
		16'hDB49: out_word = 8'h06;
		16'hDB4A: out_word = 8'h00;
		16'hDB4B: out_word = 8'hE5;
		16'hDB4C: out_word = 8'h7E;
		16'hDB4D: out_word = 8'h3F;
		16'hDB4E: out_word = 8'hF3;
		16'hDB4F: out_word = 8'h38;
		16'hDB50: out_word = 8'h07;
		16'hDB51: out_word = 8'h3E;
		16'hDB52: out_word = 8'h06;
		16'hDB53: out_word = 8'h80;
		16'hDB54: out_word = 8'hC9;
		16'hDB55: out_word = 8'h47;
		16'hDB56: out_word = 8'h23;
		16'hDB57: out_word = 8'hD8;
		16'hDB58: out_word = 8'h62;
		16'hDB59: out_word = 8'hF8;
		16'hDB5A: out_word = 8'h90;
		16'hDB5B: out_word = 8'hCB;
		16'hDB5C: out_word = 8'h3F;
		16'hDB5D: out_word = 8'h3D;
		16'hDB5E: out_word = 8'hC6;
		16'hDB5F: out_word = 8'h5F;
		16'hDB60: out_word = 8'h32;
		16'hDB61: out_word = 8'h04;
		16'hDB62: out_word = 8'h7E;
		16'hDB63: out_word = 8'hE1;
		16'hDB64: out_word = 8'hC9;
		16'hDB65: out_word = 8'hF3;
		16'hDB66: out_word = 8'hFE;
		16'hDB67: out_word = 8'h09;
		16'hDB68: out_word = 8'h20;
		16'hDB69: out_word = 8'h0F;
		16'hDB6A: out_word = 8'hCE;
		16'hDB6B: out_word = 8'h47;
		16'hDB6C: out_word = 8'hC6;
		16'hDB6D: out_word = 8'h87;
		16'hDB6E: out_word = 8'h80;
		16'hDB6F: out_word = 8'h12;
		16'hDB70: out_word = 8'h3A;
		16'hDB71: out_word = 8'h42;
		16'hDB72: out_word = 8'hF0;
		16'hDB73: out_word = 8'h43;
		16'hDB74: out_word = 8'hEC;
		16'hDB75: out_word = 8'hED;
		16'hDB76: out_word = 8'h0D;
		16'hDB77: out_word = 8'hEE;
		16'hDB78: out_word = 8'h20;
		16'hDB79: out_word = 8'h0E;
		16'hDB7A: out_word = 8'h3E;
		16'hDB7B: out_word = 8'h62;
		16'hDB7C: out_word = 8'hE2;
		16'hDB7D: out_word = 8'h3A;
		16'hDB7E: out_word = 8'h03;
		16'hDB7F: out_word = 8'h90;
		16'hDB80: out_word = 8'hA1;
		16'hDB81: out_word = 8'h03;
		16'hDB82: out_word = 8'h4E;
		16'hDB83: out_word = 8'hEE;
		16'hDB84: out_word = 8'h14;
		16'hDB85: out_word = 8'h20;
		16'hDB86: out_word = 8'h0B;
		16'hDB87: out_word = 8'h8A;
		16'hDB88: out_word = 8'hA9;
		16'hDB89: out_word = 8'h98;
		16'hDB8A: out_word = 8'h37;
		16'hDB8B: out_word = 8'hFC;
		16'hDB8C: out_word = 8'h32;
		16'hDB8D: out_word = 8'hA9;
		16'hDB8E: out_word = 8'hF1;
		16'hDB8F: out_word = 8'h16;
		16'hDB90: out_word = 8'hD7;
		16'hDB91: out_word = 8'h20;
		16'hDB92: out_word = 8'h09;
		16'hDB93: out_word = 8'h46;
		16'hDB94: out_word = 8'hD7;
		16'hDB95: out_word = 8'h5D;
		16'hDB96: out_word = 8'h7F;
		16'hDB97: out_word = 8'h4E;
		16'hDB98: out_word = 8'hF3;
		16'hDB99: out_word = 8'h17;
		16'hDB9A: out_word = 8'h20;
		16'hDB9B: out_word = 8'h06;
		16'hDB9C: out_word = 8'h74;
		16'hDB9D: out_word = 8'hE4;
		16'hDB9E: out_word = 8'h32;
		16'hDB9F: out_word = 8'h6A;
		16'hDBA0: out_word = 8'hF6;
		16'hDBA1: out_word = 8'h94;
		16'hDBA2: out_word = 8'h08;
		16'hDBA3: out_word = 8'hE9;
		16'hDBA4: out_word = 8'hBC;
		16'hDBA5: out_word = 8'hDE;
		16'hDBA6: out_word = 8'h86;
		16'hDBA7: out_word = 8'h23;
		16'hDBA8: out_word = 8'hBB;
		16'hDBA9: out_word = 8'hF8;
		16'hDBAA: out_word = 8'h01;
		16'hDBAB: out_word = 8'hC0;
		16'hDBAC: out_word = 8'hDD;
		16'hDBAD: out_word = 8'h56;
		16'hDBAE: out_word = 8'h00;
		16'hDBAF: out_word = 8'hB0;
		16'hDBB0: out_word = 8'h5E;
		16'hDBB1: out_word = 8'h6B;
		16'hDBB2: out_word = 8'hEB;
		16'hDBB3: out_word = 8'hF9;
		16'hDBB4: out_word = 8'hC9;
		16'hDBB5: out_word = 8'h24;
		16'hDBB6: out_word = 8'h22;
		16'hDBB7: out_word = 8'hD7;
		16'hDBB8: out_word = 8'h01;
		16'hDBB9: out_word = 8'h59;
		16'hDBBA: out_word = 8'h64;
		16'hDBBB: out_word = 8'h63;
		16'hDBBC: out_word = 8'h8D;
		16'hDBBD: out_word = 8'h6F;
		16'hDBBE: out_word = 8'hAF;
		16'hDBBF: out_word = 8'hA6;
		16'hDBC0: out_word = 8'h67;
		16'hDBC1: out_word = 8'hEF;
		16'hDBC2: out_word = 8'h19;
		16'hDBC3: out_word = 8'hD9;
		16'hDBC4: out_word = 8'hEE;
		16'hDBC5: out_word = 8'h9D;
		16'hDBC6: out_word = 8'hCD;
		16'hDBC7: out_word = 8'h38;
		16'hDBC8: out_word = 8'hF8;
		16'hDBC9: out_word = 8'h47;
		16'hDBCA: out_word = 8'h27;
		16'hDBCB: out_word = 8'h34;
		16'hDBCC: out_word = 8'h4F;
		16'hDBCD: out_word = 8'h68;
		16'hDBCE: out_word = 8'h84;
		16'hDBCF: out_word = 8'h67;
		16'hDBD0: out_word = 8'h4D;
		16'hDBD1: out_word = 8'hDE;
		16'hDBD2: out_word = 8'h5D;
		16'hDBD3: out_word = 8'h78;
		16'hDBD4: out_word = 8'h7F;
		16'hDBD5: out_word = 8'hA2;
		16'hDBD6: out_word = 8'h42;
		16'hDBD7: out_word = 8'h19;
		16'hDBD8: out_word = 8'h1D;
		16'hDBD9: out_word = 8'h7C;
		16'hDBDA: out_word = 8'hBA;
		16'hDBDB: out_word = 8'hFC;
		16'hDBDC: out_word = 8'hBC;
		16'hDBDD: out_word = 8'h5F;
		16'hDBDE: out_word = 8'h56;
		16'hDBDF: out_word = 8'h3E;
		16'hDBE0: out_word = 8'h15;
		16'hDBE1: out_word = 8'h91;
		16'hDBE2: out_word = 8'hF8;
		16'hDBE3: out_word = 8'hFF;
		16'hDBE4: out_word = 8'h32;
		16'hDBE5: out_word = 8'h42;
		16'hDBE6: out_word = 8'h7E;
		16'hDBE7: out_word = 8'h21;
		16'hDBE8: out_word = 8'hC2;
		16'hDBE9: out_word = 8'hC7;
		16'hDBEA: out_word = 8'h09;
		16'hDBEB: out_word = 8'h3F;
		16'hDBEC: out_word = 8'h9E;
		16'hDBED: out_word = 8'h66;
		16'hDBEE: out_word = 8'h6F;
		16'hDBEF: out_word = 8'hEB;
		16'hDBF0: out_word = 8'h3E;
		16'hDBF1: out_word = 8'h08;
		16'hDBF2: out_word = 8'h1E;
		16'hDBF3: out_word = 8'hD9;
		16'hDBF4: out_word = 8'h45;
		16'hDBF5: out_word = 8'hF7;
		16'hDBF6: out_word = 8'hFF;
		16'hDBF7: out_word = 8'hEE;
		16'hDBF8: out_word = 8'h00;
		16'hDBF9: out_word = 8'h4F;
		16'hDBFA: out_word = 8'hAF;
		16'hDBFB: out_word = 8'h18;
		16'hDBFC: out_word = 8'h13;
		16'hDBFD: out_word = 8'hCB;
		16'hDBFE: out_word = 8'h39;
		16'hDBFF: out_word = 8'hB1;
		16'hDC00: out_word = 8'h1F;
		16'hDC01: out_word = 8'h07;
		16'hDC02: out_word = 8'hFD;
		16'hDC03: out_word = 8'h47;
		16'hDC04: out_word = 8'h7E;
		16'hDC05: out_word = 8'hA3;
		16'hDC06: out_word = 8'hE1;
		16'hDC07: out_word = 8'hB1;
		16'hDC08: out_word = 8'h77;
		16'hDC09: out_word = 8'h2C;
		16'hDC0A: out_word = 8'hD7;
		16'hDC0B: out_word = 8'hA2;
		16'hDC0C: out_word = 8'hFF;
		16'hDC0D: out_word = 8'hAB;
		16'hDC0E: out_word = 8'h24;
		16'hDC0F: out_word = 8'h08;
		16'hDC10: out_word = 8'h3D;
		16'hDC11: out_word = 8'hC2;
		16'hDC12: out_word = 8'h38;
		16'hDC13: out_word = 8'h7E;
		16'hDC14: out_word = 8'hFE;
		16'hDC15: out_word = 8'h1E;
		16'hDC16: out_word = 8'h00;
		16'hDC17: out_word = 8'h1C;
		16'hDC18: out_word = 8'h28;
		16'hDC19: out_word = 8'h0C;
		16'hDC1A: out_word = 8'h25;
		16'hDC1B: out_word = 8'h1D;
		16'hDC1C: out_word = 8'hDB;
		16'hDC1D: out_word = 8'hFD;
		16'hDC1E: out_word = 8'h66;
		16'hDC1F: out_word = 8'h67;
		16'hDC20: out_word = 8'h73;
		16'hDC21: out_word = 8'hD9;
		16'hDC22: out_word = 8'h5B;
		16'hDC23: out_word = 8'h1F;
		16'hDC24: out_word = 8'h03;
		16'hDC25: out_word = 8'hFF;
		16'hDC26: out_word = 8'h8D;
		16'hDC27: out_word = 8'h81;
		16'hDC28: out_word = 8'hC0;
		16'hDC29: out_word = 8'h13;
		16'hDC2A: out_word = 8'hE0;
		16'hDC2B: out_word = 8'h7F;
		16'hDC2C: out_word = 8'hFF;
		16'hDC2D: out_word = 8'hF0;
		16'hDC2E: out_word = 8'h3F;
		16'hDC2F: out_word = 8'hF8;
		16'hDC30: out_word = 8'h1F;
		16'hDC31: out_word = 8'hFC;
		16'hDC32: out_word = 8'h0F;
		16'hDC33: out_word = 8'hFE;
		16'hDC34: out_word = 8'h07;
		16'hDC35: out_word = 8'hAC;
		16'hDC36: out_word = 8'hC5;
		16'hDC37: out_word = 8'h6E;
		16'hDC38: out_word = 8'hD5;
		16'hDC39: out_word = 8'hF6;
		16'hDC3A: out_word = 8'h10;
		16'hDC3B: out_word = 8'hB3;
		16'hDC3C: out_word = 8'h1C;
		16'hDC3D: out_word = 8'hFE;
		16'hDC3E: out_word = 8'h12;
		16'hDC3F: out_word = 8'h6B;
		16'hDC40: out_word = 8'h4D;
		16'hDC41: out_word = 8'h79;
		16'hDC42: out_word = 8'h9A;
		16'hDC43: out_word = 8'hAC;
		16'hDC44: out_word = 8'h4F;
		16'hDC45: out_word = 8'h78;
		16'hDC46: out_word = 8'h7F;
		16'hDC47: out_word = 8'hFB;
		16'hDC48: out_word = 8'hCD;
		16'hDC49: out_word = 8'hB0;
		16'hDC4A: out_word = 8'h22;
		16'hDC4B: out_word = 8'hEB;
		16'hDC4C: out_word = 8'hDD;
		16'hDC4D: out_word = 8'hE5;
		16'hDC4E: out_word = 8'hE1;
		16'hDC4F: out_word = 8'h98;
		16'hDC50: out_word = 8'h23;
		16'hDC51: out_word = 8'hFF;
		16'hDC52: out_word = 8'h46;
		16'hDC53: out_word = 8'h94;
		16'hDC54: out_word = 8'h05;
		16'hDC55: out_word = 8'h1A;
		16'hDC56: out_word = 8'hFC;
		16'hDC57: out_word = 8'h77;
		16'hDC58: out_word = 8'h7F;
		16'hDC59: out_word = 8'hD5;
		16'hDC5A: out_word = 8'h48;
		16'hDC5B: out_word = 8'hCD;
		16'hDC5C: out_word = 8'h84;
		16'hDC5D: out_word = 8'h3E;
		16'hDC5E: out_word = 8'h0D;
		16'hDC5F: out_word = 8'h20;
		16'hDC60: out_word = 8'hFA;
		16'hDC61: out_word = 8'h14;
		16'hDC62: out_word = 8'h81;
		16'hDC63: out_word = 8'h2C;
		16'hDC64: out_word = 8'hD1;
		16'hDC65: out_word = 8'hD5;
		16'hDC66: out_word = 8'h38;
		16'hDC67: out_word = 8'h12;
		16'hDC68: out_word = 8'h60;
		16'hDC69: out_word = 8'h40;
		16'hDC6A: out_word = 8'hA3;
		16'hDC6B: out_word = 8'hAE;
		16'hDC6C: out_word = 8'h23;
		16'hDC6D: out_word = 8'h53;
		16'hDC6E: out_word = 8'h9D;
		16'hDC6F: out_word = 8'hC5;
		16'hDC70: out_word = 8'hEA;
		16'hDC71: out_word = 8'h10;
		16'hDC72: out_word = 8'hFB;
		16'hDC73: out_word = 8'hB9;
		16'hDC74: out_word = 8'hC1;
		16'hDC75: out_word = 8'hC7;
		16'hDC76: out_word = 8'hC6;
		16'hDC77: out_word = 8'hDC;
		16'hDC78: out_word = 8'h0E;
		16'hDC79: out_word = 8'h57;
		16'hDC7A: out_word = 8'hC5;
		16'hDC7B: out_word = 8'h07;
		16'hDC7C: out_word = 8'h0D;
		16'hDC7D: out_word = 8'h5F;
		16'hDC7E: out_word = 8'hFF;
		16'hDC7F: out_word = 8'hE1;
		16'hDC80: out_word = 8'h24;
		16'hDC81: out_word = 8'h0E;
		16'hDC82: out_word = 8'h40;
		16'hDC83: out_word = 8'hC5;
		16'hDC84: out_word = 8'hE5;
		16'hDC85: out_word = 8'h43;
		16'hDC86: out_word = 8'hCD;
		16'hDC87: out_word = 8'hE2;
		16'hDC88: out_word = 8'hFB;
		16'hDC89: out_word = 8'h7E;
		16'hDC8A: out_word = 8'h42;
		16'hDC8B: out_word = 8'h7B;
		16'hDC8C: out_word = 8'h0C;
		16'hDC8D: out_word = 8'h7F;
		16'hDC8E: out_word = 8'hE1;
		16'hDC8F: out_word = 8'hC1;
		16'hDC90: out_word = 8'h9F;
		16'hDC91: out_word = 8'hFA;
		16'hDC92: out_word = 8'h43;
		16'hDC93: out_word = 8'h7E;
		16'hDC94: out_word = 8'hB1;
		16'hDC95: out_word = 8'hCB;
		16'hDC96: out_word = 8'h09;
		16'hDC97: out_word = 8'hD3;
		16'hDC98: out_word = 8'h30;
		16'hDC99: out_word = 8'h03;
		16'hDC9A: out_word = 8'h5B;
		16'hDC9B: out_word = 8'h10;
		16'hDC9C: out_word = 8'hF6;
		16'hDC9D: out_word = 8'h3E;
		16'hDC9E: out_word = 8'h55;
		16'hDC9F: out_word = 8'hC9;
		16'hDCA0: out_word = 8'hCD;
		16'hDCA1: out_word = 8'h2E;
		16'hDCA2: out_word = 8'h7D;
		16'hDCA3: out_word = 8'h41;
		16'hDCA4: out_word = 8'hEF;
		16'hDCA5: out_word = 8'hFF;
		16'hDCA6: out_word = 8'h10;
		16'hDCA7: out_word = 8'hF8;
		16'hDCA8: out_word = 8'hC9;
		16'hDCA9: out_word = 8'h7B;
		16'hDCAA: out_word = 8'hC6;
		16'hDCAB: out_word = 8'h20;
		16'hDCAC: out_word = 8'h5F;
		16'hDCAD: out_word = 8'hD0;
		16'hDCAE: out_word = 8'h87;
		16'hDCAF: out_word = 8'h7A;
		16'hDCB0: out_word = 8'h08;
		16'hDCB1: out_word = 8'hAA;
		16'hDCB2: out_word = 8'h57;
		16'hDCB3: out_word = 8'h64;
		16'hDCB4: out_word = 8'hDB;
		16'hDCB5: out_word = 8'hD5;
		16'hDCB6: out_word = 8'hE5;
		16'hDCB7: out_word = 8'h13;
		16'hDCB8: out_word = 8'h9D;
		16'hDCB9: out_word = 8'hE7;
		16'hDCBA: out_word = 8'hCF;
		16'hDCBB: out_word = 8'hD1;
		16'hDCBC: out_word = 8'h23;
		16'hDCBD: out_word = 8'h3C;
		16'hDCBE: out_word = 8'h9F;
		16'hDCBF: out_word = 8'h10;
		16'hDCC0: out_word = 8'hEF;
		16'hDCC1: out_word = 8'hC9;
		16'hDCC2: out_word = 8'h7C;
		16'hDCC3: out_word = 8'h18;
		16'hDCC4: out_word = 8'h33;
		16'hDCC5: out_word = 8'h3A;
		16'hDCC6: out_word = 8'h7D;
		16'hDCC7: out_word = 8'hF5;
		16'hDCC8: out_word = 8'h0B;
		16'hDCC9: out_word = 8'h3D;
		16'hDCCA: out_word = 8'hCD;
		16'hDCCB: out_word = 8'hF3;
		16'hDCCC: out_word = 8'h3C;
		16'hDCCD: out_word = 8'h7F;
		16'hDCCE: out_word = 8'hF1;
		16'hDCCF: out_word = 8'hE6;
		16'hDCD0: out_word = 8'h4E;
		16'hDCD1: out_word = 8'h0A;
		16'hDCD2: out_word = 8'hF0;
		16'hDCD3: out_word = 8'h3F;
		16'hDCD4: out_word = 8'hCE;
		16'hDCD5: out_word = 8'h30;
		16'hDCD6: out_word = 8'h27;
		16'hDCD7: out_word = 8'h20;
		16'hDCD8: out_word = 8'h7F;
		16'hDCD9: out_word = 8'h42;
		16'hDCDA: out_word = 8'h20;
		16'hDCDB: out_word = 8'h89;
		16'hDCDC: out_word = 8'h06;
		16'hDCDD: out_word = 8'h80;
		16'hDCDE: out_word = 8'hF9;
		16'hDCDF: out_word = 8'h38;
		16'hDCE0: out_word = 8'h02;
		16'hDCE1: out_word = 8'h3E;
		16'hDCE2: out_word = 8'h2E;
		16'hDCE3: out_word = 8'hD5;
		16'hDCE4: out_word = 8'h99;
		16'hDCE5: out_word = 8'hF8;
		16'hDCE6: out_word = 8'h87;
		16'hDCE7: out_word = 8'h6F;
		16'hDCE8: out_word = 8'h26;
		16'hDCE9: out_word = 8'h0F;
		16'hDCEA: out_word = 8'h29;
		16'hDCEB: out_word = 8'hFC;
		16'hDCEC: out_word = 8'h06;
		16'hDCED: out_word = 8'h04;
		16'hDCEE: out_word = 8'h7E;
		16'hDCEF: out_word = 8'h2F;
		16'hDCF0: out_word = 8'hB6;
		16'hDCF1: out_word = 8'h2C;
		16'hDCF2: out_word = 8'hEB;
		16'hDCF3: out_word = 8'h77;
		16'hDCF4: out_word = 8'h8A;
		16'hDCF5: out_word = 8'h24;
		16'hDCF6: out_word = 8'hD9;
		16'hDCF7: out_word = 8'hF8;
		16'hDCF8: out_word = 8'h10;
		16'hDCF9: out_word = 8'h9A;
		16'hDCFA: out_word = 8'hEE;
		16'hDCFB: out_word = 8'h87;
		16'hDCFC: out_word = 8'h7A;
		16'hDCFD: out_word = 8'h7F;
		16'hDCFE: out_word = 8'hC5;
		16'hDCFF: out_word = 8'hC6;
		16'hDD00: out_word = 8'h4F;
		16'hDD01: out_word = 8'h57;
		16'hDD02: out_word = 8'h3E;
		16'hDD03: out_word = 8'h07;
		16'hDD04: out_word = 8'h12;
		16'hDD05: out_word = 8'hD1;
		16'hDD06: out_word = 8'hDE;
		16'hDD07: out_word = 8'h1C;
		16'hDD08: out_word = 8'hC0;
		16'hDD09: out_word = 8'h9B;
		16'hDD0A: out_word = 8'h43;
		16'hDD0B: out_word = 8'h51;
		16'hDD0C: out_word = 8'hCC;
		16'hDD0D: out_word = 8'hAF;
		16'hDD0E: out_word = 8'hD9;
		16'hDD0F: out_word = 8'h12;
		16'hDD10: out_word = 8'h14;
		16'hDD11: out_word = 8'h8D;
		16'hDD12: out_word = 8'hFE;
		16'hDD13: out_word = 8'h18;
		16'hDD14: out_word = 8'hD5;
		16'hDD15: out_word = 8'h16;
		16'hDD16: out_word = 8'h29;
		16'hDD17: out_word = 8'h93;
		16'hDD18: out_word = 8'hB0;
		16'hDD19: out_word = 8'h89;
		16'hDD1A: out_word = 8'h0C;
		16'hDD1B: out_word = 8'hED;
		16'hDD1C: out_word = 8'hC3;
		16'hDD1D: out_word = 8'h53;
		16'hDD1E: out_word = 8'h9D;
		16'hDD1F: out_word = 8'h4F;
		16'hDD20: out_word = 8'hF2;
		16'hDD21: out_word = 8'h7E;
		16'hDD22: out_word = 8'hFE;
		16'hDD23: out_word = 8'hFF;
		16'hDD24: out_word = 8'hC8;
		16'hDD25: out_word = 8'h06;
		16'hDD26: out_word = 8'h44;
		16'hDD27: out_word = 8'h0C;
		16'hDD28: out_word = 8'hCB;
		16'hDD29: out_word = 8'hFF;
		16'hDD2A: out_word = 8'h6A;
		16'hDD2B: out_word = 8'h28;
		16'hDD2C: out_word = 8'hF4;
		16'hDD2D: out_word = 8'h18;
		16'hDD2E: out_word = 8'hE1;
		16'hDD2F: out_word = 8'hE5;
		16'hDD30: out_word = 8'h7A;
		16'hDD31: out_word = 8'hCD;
		16'hDD32: out_word = 8'hFE;
		16'hDD33: out_word = 8'h9E;
		16'hDD34: out_word = 8'h0E;
		16'hDD35: out_word = 8'h7B;
		16'hDD36: out_word = 8'h85;
		16'hDD37: out_word = 8'h6F;
		16'hDD38: out_word = 8'hEB;
		16'hDD39: out_word = 8'hE1;
		16'hDD3A: out_word = 8'h5A;
		16'hDD3B: out_word = 8'hF0;
		16'hDD3C: out_word = 8'h3E;
		16'hDD3D: out_word = 8'hE7;
		16'hDD3E: out_word = 8'h18;
		16'hDD3F: out_word = 8'hF6;
		16'hDD40: out_word = 8'hED;
		16'hDD41: out_word = 8'h5B;
		16'hDD42: out_word = 8'hE3;
		16'hDD43: out_word = 8'h17;
		16'hDD44: out_word = 8'h21;
		16'hDD45: out_word = 8'h90;
		16'hDD46: out_word = 8'hF7;
		16'hDD47: out_word = 8'hFF;
		16'hDD48: out_word = 8'hDD;
		16'hDD49: out_word = 8'h4E;
		16'hDD4A: out_word = 8'h03;
		16'hDD4B: out_word = 8'hFD;
		16'hDD4C: out_word = 8'hCB;
		16'hDD4D: out_word = 8'h37;
		16'hDD4E: out_word = 8'h56;
		16'hDD4F: out_word = 8'h28;
		16'hDD50: out_word = 8'hEE;
		16'hDD51: out_word = 8'h01;
		16'hDD52: out_word = 8'h0D;
		16'hDD53: out_word = 8'h06;
		16'hDD54: out_word = 8'hBA;
		16'hDD55: out_word = 8'hD4;
		16'hDD56: out_word = 8'h34;
		16'hDD57: out_word = 8'hBA;
		16'hDD58: out_word = 8'h38;
		16'hDD59: out_word = 8'hEB;
		16'hDD5A: out_word = 8'hF2;
		16'hDD5B: out_word = 8'h09;
		16'hDD5C: out_word = 8'h73;
		16'hDD5D: out_word = 8'hAE;
		16'hDD5E: out_word = 8'h47;
		16'hDD5F: out_word = 8'h2E;
		16'hDD60: out_word = 8'h19;
		16'hDD61: out_word = 8'h9B;
		16'hDD62: out_word = 8'hF3;
		16'hDD63: out_word = 8'hC5;
		16'hDD64: out_word = 8'h2C;
		16'hDD65: out_word = 8'hBB;
		16'hDD66: out_word = 8'hF0;
		16'hDD67: out_word = 8'h22;
		16'hDD68: out_word = 8'h94;
		16'hDD69: out_word = 8'hE3;
		16'hDD6A: out_word = 8'h99;
		16'hDD6B: out_word = 8'hE2;
		16'hDD6C: out_word = 8'h5A;
		16'hDD6D: out_word = 8'hD3;
		16'hDD6E: out_word = 8'hFF;
		16'hDD6F: out_word = 8'h4E;
		16'hDD70: out_word = 8'h05;
		16'hDD71: out_word = 8'h7E;
		16'hDD72: out_word = 8'h12;
		16'hDD73: out_word = 8'h71;
		16'hDD74: out_word = 8'h2C;
		16'hDD75: out_word = 8'h1C;
		16'hDD76: out_word = 8'h10;
		16'hDD77: out_word = 8'hAF;
		16'hDD78: out_word = 8'hF9;
		16'hDD79: out_word = 8'h5C;
		16'hDD7A: out_word = 8'hE1;
		16'hDD7B: out_word = 8'hEB;
		16'hDD7C: out_word = 8'hE5;
		16'hDD7D: out_word = 8'h53;
		16'hDD7E: out_word = 8'h47;
		16'hDD7F: out_word = 8'hB4;
		16'hDD80: out_word = 8'hF8;
		16'hDD81: out_word = 8'hD6;
		16'hDD82: out_word = 8'hFE;
		16'hDD83: out_word = 8'h09;
		16'hDD84: out_word = 8'hC1;
		16'hDD85: out_word = 8'h76;
		16'hDD86: out_word = 8'hE5;
		16'hDD87: out_word = 8'h2C;
		16'hDD88: out_word = 8'h14;
		16'hDD89: out_word = 8'h34;
		16'hDD8A: out_word = 8'hFC;
		16'hDD8B: out_word = 8'hC1;
		16'hDD8C: out_word = 8'hD1;
		16'hDD8D: out_word = 8'hE1;
		16'hDD8E: out_word = 8'h6C;
		16'hDD8F: out_word = 8'hC9;
		16'hDD90: out_word = 8'h68;
		16'hDD91: out_word = 8'h01;
		16'hDD92: out_word = 8'h44;
		16'hDD93: out_word = 8'h0B;
		16'hDD94: out_word = 8'hE9;
		16'hDD95: out_word = 8'h61;
		16'hDD96: out_word = 8'h39;
		16'hDD97: out_word = 8'hFA;
		16'hDD98: out_word = 8'hE3;
		16'hDD99: out_word = 8'hBF;
		16'hDD9A: out_word = 8'h7D;
		16'hDD9B: out_word = 8'h12;
		16'hDD9C: out_word = 8'h3F;
		16'hDD9D: out_word = 8'h77;
		16'hDD9E: out_word = 8'h13;
		16'hDD9F: out_word = 8'h78;
		16'hDDA0: out_word = 8'hB1;
		16'hDDA1: out_word = 8'hC8;
		16'hDDA2: out_word = 8'h0B;
		16'hDDA3: out_word = 8'h06;
		16'hDDA4: out_word = 8'h71;
		16'hDDA5: out_word = 8'h74;
		16'hDDA6: out_word = 8'hF6;
		16'hDDA7: out_word = 8'h70;
		16'hDDA8: out_word = 8'h13;
		16'hDDA9: out_word = 8'h53;
		16'hDDAA: out_word = 8'hE1;
		16'hDDAB: out_word = 8'hA7;
		16'hDDAC: out_word = 8'h28;
		16'hDDAD: out_word = 8'h06;
		16'hDDAE: out_word = 8'h42;
		16'hDDAF: out_word = 8'h35;
		16'hDDB0: out_word = 8'hFC;
		16'hDDB1: out_word = 8'hC3;
		16'hDDB2: out_word = 8'hE2;
		16'hDDB3: out_word = 8'h7F;
		16'hDDB4: out_word = 8'hCD;
		16'hDDB5: out_word = 8'h94;
		16'hDDB6: out_word = 8'h63;
		16'hDDB7: out_word = 8'h5D;
		16'hDDB8: out_word = 8'hE6;
		16'hDDB9: out_word = 8'h7B;
		16'hDDBA: out_word = 8'h7A;
		16'hDDBB: out_word = 8'h3A;
		16'hDDBC: out_word = 8'h1C;
		16'hDDBD: out_word = 8'hBD;
		16'hDDBE: out_word = 8'h33;
		16'hDDBF: out_word = 8'h14;
		16'hDDC0: out_word = 8'h1F;
		16'hDDC1: out_word = 8'h21;
		16'hDDC2: out_word = 8'h55;
		16'hDDC3: out_word = 8'hE6;
		16'hDDC4: out_word = 8'h6C;
		16'hDDC5: out_word = 8'hCB;
		16'hDDC6: out_word = 8'h5E;
		16'hDDC7: out_word = 8'h3A;
		16'hDDC8: out_word = 8'h12;
		16'hDDC9: out_word = 8'h67;
		16'hDDCA: out_word = 8'h34;
		16'hDDCB: out_word = 8'h13;
		16'hDDCC: out_word = 8'h5A;
		16'hDDCD: out_word = 8'hC0;
		16'hDDCE: out_word = 8'h20;
		16'hDDCF: out_word = 8'hDC;
		16'hDDD0: out_word = 8'h11;
		16'hDDD1: out_word = 8'h29;
		16'hDDD2: out_word = 8'h5A;
		16'hDDD3: out_word = 8'hFE;
		16'hDDD4: out_word = 8'h06;
		16'hDDD5: out_word = 8'h08;
		16'hDDD6: out_word = 8'h7E;
		16'hDDD7: out_word = 8'h23;
		16'hDDD8: out_word = 8'hCD;
		16'hDDD9: out_word = 8'h4B;
		16'hDDDA: out_word = 8'h80;
		16'hDDDB: out_word = 8'h79;
		16'hDDDC: out_word = 8'h3E;
		16'hDDDD: out_word = 8'hC3;
		16'hDDDE: out_word = 8'h5E;
		16'hDDDF: out_word = 8'h64;
		16'hDDE0: out_word = 8'hF2;
		16'hDDE1: out_word = 8'h58;
		16'hDDE2: out_word = 8'hC4;
		16'hDDE3: out_word = 8'hD4;
		16'hDDE4: out_word = 8'hD5;
		16'hDDE5: out_word = 8'h3E;
		16'hDDE6: out_word = 8'h6E;
		16'hDDE7: out_word = 8'hC6;
		16'hDDE8: out_word = 8'h90;
		16'hDDE9: out_word = 8'h47;
		16'hDDEA: out_word = 8'hFC;
		16'hDDEB: out_word = 8'h01;
		16'hDDEC: out_word = 8'hFF;
		16'hDDED: out_word = 8'h0B;
		16'hDDEE: out_word = 8'h00;
		16'hDDEF: out_word = 8'h09;
		16'hDDF0: out_word = 8'h7E;
		16'hDDF1: out_word = 8'hED;
		16'hDDF2: out_word = 8'h42;
		16'hDDF3: out_word = 8'hE6;
		16'hDDF4: out_word = 8'h10;
		16'hDDF5: out_word = 8'h81;
		16'hDDF6: out_word = 8'h3E;
		16'hDDF7: out_word = 8'h20;
		16'hDDF8: out_word = 8'h89;
		16'hDDF9: out_word = 8'h02;
		16'hDDFA: out_word = 8'h01;
		16'hDDFB: out_word = 8'hFD;
		16'hDDFC: out_word = 8'hD1;
		16'hDDFD: out_word = 8'hCD;
		16'hDDFE: out_word = 8'h14;
		16'hDDFF: out_word = 8'h80;
		16'hDE00: out_word = 8'h18;
		16'hDE01: out_word = 8'hCF;
		16'hDE02: out_word = 8'hA0;
		16'hDE03: out_word = 8'h8F;
		16'hDE04: out_word = 8'hD6;
		16'hDE05: out_word = 8'hB9;
		16'hDE06: out_word = 8'h10;
		16'hDE07: out_word = 8'hFC;
		16'hDE08: out_word = 8'hC7;
		16'hDE09: out_word = 8'h7C;
		16'hDE0A: out_word = 8'hB5;
		16'hDE0B: out_word = 8'hC8;
		16'hDE0C: out_word = 8'h37;
		16'hDE0D: out_word = 8'h89;
		16'hDE0E: out_word = 8'hE0;
		16'hDE0F: out_word = 8'h03;
		16'hDE10: out_word = 8'h6C;
		16'hDE11: out_word = 8'h85;
		16'hDE12: out_word = 8'hCE;
		16'hDE13: out_word = 8'h02;
		16'hDE14: out_word = 8'hD6;
		16'hDE15: out_word = 8'hF5;
		16'hDE16: out_word = 8'hBE;
		16'hDE17: out_word = 8'h0F;
		16'hDE18: out_word = 8'h96;
		16'hDE19: out_word = 8'h81;
		16'hDE1A: out_word = 8'h34;
		16'hDE1B: out_word = 8'hCD;
		16'hDE1C: out_word = 8'h81;
		16'hDE1D: out_word = 8'hBE;
		16'hDE1E: out_word = 8'h7B;
		16'hDE1F: out_word = 8'hF9;
		16'hDE20: out_word = 8'hE9;
		16'hDE21: out_word = 8'h23;
		16'hDE22: out_word = 8'hE7;
		16'hDE23: out_word = 8'h79;
		16'hDE24: out_word = 8'h5F;
		16'hDE25: out_word = 8'hC3;
		16'hDE26: out_word = 8'hB2;
		16'hDE27: out_word = 8'h80;
		16'hDE28: out_word = 8'h75;
		16'hDE29: out_word = 8'hAD;
		16'hDE2A: out_word = 8'h10;
		16'hDE2B: out_word = 8'hBC;
		16'hDE2C: out_word = 8'hC6;
		16'hDE2D: out_word = 8'h7D;
		16'hDE2E: out_word = 8'hD1;
		16'hDE2F: out_word = 8'hD2;
		16'hDE30: out_word = 8'h4F;
		16'hDE31: out_word = 8'hF5;
		16'hDE32: out_word = 8'h06;
		16'hDE33: out_word = 8'h00;
		16'hDE34: out_word = 8'h7A;
		16'hDE35: out_word = 8'hB3;
		16'hDE36: out_word = 8'h7F;
		16'hDE37: out_word = 8'hC6;
		16'hDE38: out_word = 8'h39;
		16'hDE39: out_word = 8'h81;
		16'hDE3A: out_word = 8'hC8;
		16'hDE3B: out_word = 8'hAF;
		16'hDE3C: out_word = 8'h3F;
		16'hDE3D: out_word = 8'hB7;
		16'hDE3E: out_word = 8'hEB;
		16'hDE3F: out_word = 8'h30;
		16'hDE40: out_word = 8'h1F;
		16'hDE41: out_word = 8'h57;
		16'hDE42: out_word = 8'h5F;
		16'hDE43: out_word = 8'hDC;
		16'hDE44: out_word = 8'h18;
		16'hDE45: out_word = 8'h1B;
		16'hDE46: out_word = 8'hF2;
		16'hDE47: out_word = 8'hCC;
		16'hDE48: out_word = 8'hEB;
		16'hDE49: out_word = 8'hA7;
		16'hDE4A: out_word = 8'hF1;
		16'hDE4B: out_word = 8'h09;
		16'hDE4C: out_word = 8'hFC;
		16'hDE4D: out_word = 8'hF0;
		16'hDE4E: out_word = 8'h04;
		16'hDE4F: out_word = 8'h1B;
		16'hDE50: out_word = 8'h7B;
		16'hDE51: out_word = 8'h18;
		16'hDE52: out_word = 8'h0B;
		16'hDE53: out_word = 8'hFE;
		16'hDE54: out_word = 8'hF8;
		16'hDE55: out_word = 8'hED;
		16'hDE56: out_word = 8'h52;
		16'hDE57: out_word = 8'h19;
		16'hDE58: out_word = 8'h28;
		16'hDE59: out_word = 8'h02;
		16'hDE5A: out_word = 8'h30;
		16'hDE5B: out_word = 8'h30;
		16'hDE5C: out_word = 8'h1E;
		16'hDE5D: out_word = 8'h1B;
		16'hDE5E: out_word = 8'hDD;
		16'hDE5F: out_word = 8'h77;
		16'hDE60: out_word = 8'h0F;
		16'hDE61: out_word = 8'h2C;
		16'hDE62: out_word = 8'h73;
		16'hDE63: out_word = 8'hEE;
		16'hDE64: out_word = 8'hC2;
		16'hDE65: out_word = 8'h72;
		16'hDE66: out_word = 8'h13;
		16'hDE67: out_word = 8'h68;
		16'hDE68: out_word = 8'hA4;
		16'hDE69: out_word = 8'h86;
		16'hDE6A: out_word = 8'h84;
		16'hDE6B: out_word = 8'h4C;
		16'hDE6C: out_word = 8'hD3;
		16'hDE6D: out_word = 8'h87;
		16'hDE6E: out_word = 8'h56;
		16'hDE6F: out_word = 8'hA1;
		16'hDE70: out_word = 8'h67;
		16'hDE71: out_word = 8'h2E;
		16'hDE72: out_word = 8'h01;
		16'hDE73: out_word = 8'h7D;
		16'hDE74: out_word = 8'hB7;
		16'hDE75: out_word = 8'hDB;
		16'hDE76: out_word = 8'h4E;
		16'hDE77: out_word = 8'h5E;
		16'hDE78: out_word = 8'h42;
		16'hDE79: out_word = 8'h3E;
		16'hDE7A: out_word = 8'hF1;
		16'hDE7B: out_word = 8'h47;
		16'hDE7C: out_word = 8'h24;
		16'hDE7D: out_word = 8'h36;
		16'hDE7E: out_word = 8'h01;
		16'hDE7F: out_word = 8'hBC;
		16'hDE80: out_word = 8'h62;
		16'hDE81: out_word = 8'h7F;
		16'hDE82: out_word = 8'h29;
		16'hDE83: out_word = 8'h7C;
		16'hDE84: out_word = 8'hD6;
		16'hDE85: out_word = 8'h07;
		16'hDE86: out_word = 8'h67;
		16'hDE87: out_word = 8'h2C;
		16'hDE88: out_word = 8'h11;
		16'hDE89: out_word = 8'hFE;
		16'hDE8A: out_word = 8'hC8;
		16'hDE8B: out_word = 8'hF8;
		16'hDE8C: out_word = 8'h1A;
		16'hDE8D: out_word = 8'h2F;
		16'hDE8E: out_word = 8'h77;
		16'hDE8F: out_word = 8'h24;
		16'hDE90: out_word = 8'h1C;
		16'hDE91: out_word = 8'hC7;
		16'hDE92: out_word = 8'h13;
		16'hDE93: out_word = 8'hFB;
		16'hDE94: out_word = 8'hE1;
		16'hDE95: out_word = 8'hD8;
		16'hDE96: out_word = 8'hC1;
		16'hDE97: out_word = 8'h82;
		16'hDE98: out_word = 8'hF8;
		16'hDE99: out_word = 8'h96;
		16'hDE9A: out_word = 8'hF5;
		16'hDE9B: out_word = 8'h1C;
		16'hDE9C: out_word = 8'h38;
		16'hDE9D: out_word = 8'hFB;
		16'hDE9E: out_word = 8'hFF;
		16'hDE9F: out_word = 8'hC9;
		16'hDEA0: out_word = 8'hF3;
		16'hDEA1: out_word = 8'hC5;
		16'hDEA2: out_word = 8'h01;
		16'hDEA3: out_word = 8'hF7;
		16'hDEA4: out_word = 8'hEF;
		16'hDEA5: out_word = 8'h3E;
		16'hDEA6: out_word = 8'h80;
		16'hDEA7: out_word = 8'hF1;
		16'hDEA8: out_word = 8'hED;
		16'hDEA9: out_word = 8'h79;
		16'hDEAA: out_word = 8'h06;
		16'hDEAB: out_word = 8'hDF;
		16'hDEAC: out_word = 8'h22;
		16'hDEAD: out_word = 8'h61;
		16'hDEAE: out_word = 8'h40;
		16'hDEAF: out_word = 8'hBF;
		16'hDEB0: out_word = 8'hEC;
		16'hDEB1: out_word = 8'h68;
		16'hDEB2: out_word = 8'h18;
		16'hDEB3: out_word = 8'h11;
		16'hDEB4: out_word = 8'hE7;
		16'hDEB5: out_word = 8'hED;
		16'hDEB6: out_word = 8'h69;
		16'hDEB7: out_word = 8'h3E;
		16'hDEB8: out_word = 8'h00;
		16'hDEB9: out_word = 8'h0A;
		16'hDEBA: out_word = 8'hEF;
		16'hDEBB: out_word = 8'hBB;
		16'hDEBC: out_word = 8'h6C;
		16'hDEBD: out_word = 8'h7D;
		16'hDEBE: out_word = 8'hFF;
		16'hDEBF: out_word = 8'hA7;
		16'hDEC0: out_word = 8'hC9;
		16'hDEC1: out_word = 8'h4D;
		16'hDEC2: out_word = 8'h26;
		16'hDEC3: out_word = 8'hF0;
		16'hDEC4: out_word = 8'hCD;
		16'hDEC5: out_word = 8'h13;
		16'hDEC6: out_word = 8'h82;
		16'hDEC7: out_word = 8'h16;
		16'hDEC8: out_word = 8'h00;
		16'hDEC9: out_word = 8'h2F;
		16'hDECA: out_word = 8'hB9;
		16'hDECB: out_word = 8'hC8;
		16'hDECC: out_word = 8'h3C;
		16'hDECD: out_word = 8'h1B;
		16'hDECE: out_word = 8'hF3;
		16'hDECF: out_word = 8'h3D;
		16'hDED0: out_word = 8'hFD;
		16'hDED1: out_word = 8'hD5;
		16'hDED2: out_word = 8'h12;
		16'hDED3: out_word = 8'h13;
		16'hDED4: out_word = 8'h06;
		16'hDED5: out_word = 8'h0F;
		16'hDED6: out_word = 8'h24;
		16'hDED7: out_word = 8'h0F;
		16'hDED8: out_word = 8'hF1;
		16'hDED9: out_word = 8'hF8;
		16'hDEDA: out_word = 8'h10;
		16'hDEDB: out_word = 8'hF8;
		16'hDEDC: out_word = 8'hD1;
		16'hDEDD: out_word = 8'hFA;
		16'hDEDE: out_word = 8'h62;
		16'hDEDF: out_word = 8'h6B;
		16'hDEE0: out_word = 8'h06;
		16'hDEE1: out_word = 8'h0C;
		16'hDEE2: out_word = 8'h1A;
		16'hDEE3: out_word = 8'h84;
		16'hDEE4: out_word = 8'h17;
		16'hDEE5: out_word = 8'h13;
		16'hDEE6: out_word = 8'hF7;
		16'hDEE7: out_word = 8'h56;
		16'hDEE8: out_word = 8'h01;
		16'hDEE9: out_word = 8'h0C;
		16'hDEEA: out_word = 8'h00;
		16'hDEEB: out_word = 8'h7F;
		16'hDEEC: out_word = 8'h80;
		16'hDEED: out_word = 8'hEB;
		16'hDEEE: out_word = 8'h36;
		16'hDEEF: out_word = 8'h87;
		16'hDEF0: out_word = 8'h20;
		16'hDEF1: out_word = 8'h79;
		16'hDEF2: out_word = 8'hFB;
		16'hDEF3: out_word = 8'hE6;
		16'hDEF4: out_word = 8'h1F;
		16'hDEF5: out_word = 8'hCD;
		16'hDEF6: out_word = 8'h09;
		16'hDEF7: out_word = 8'h83;
		16'hDEF8: out_word = 8'hAF;
		16'hDEF9: out_word = 8'h8F;
		16'hDEFA: out_word = 8'h79;
		16'hDEFB: out_word = 8'hBB;
		16'hDEFC: out_word = 8'h0F;
		16'hDEFD: out_word = 8'hA1;
		16'hDEFE: out_word = 8'h04;
		16'hDEFF: out_word = 8'hF4;
		16'hDF00: out_word = 8'h36;
		16'hDF01: out_word = 8'h2E;
		16'hDF02: out_word = 8'h23;
		16'hDF03: out_word = 8'hEF;
		16'hDF04: out_word = 8'h41;
		16'hDF05: out_word = 8'hFA;
		16'hDF06: out_word = 8'h66;
		16'hDF07: out_word = 8'h32;
		16'hDF08: out_word = 8'hFD;
		16'hDF09: out_word = 8'h30;
		16'hDF0A: out_word = 8'h17;
		16'hDF0B: out_word = 8'h78;
		16'hDF0C: out_word = 8'hE6;
		16'hDF0D: out_word = 8'h3F;
		16'hDF0E: out_word = 8'h73;
		16'hDF0F: out_word = 8'hE0;
		16'hDF10: out_word = 8'h70;
		16'hDF11: out_word = 8'hC0;
		16'hDF12: out_word = 8'hFD;
		16'hDF13: out_word = 8'hEB;
		16'hDF14: out_word = 8'h21;
		16'hDF15: out_word = 8'h42;
		16'hDF16: out_word = 8'h6C;
		16'hDF17: out_word = 8'h01;
		16'hDF18: out_word = 8'h05;
		16'hDF19: out_word = 8'h7B;
		16'hDF1A: out_word = 8'h5C;
		16'hDF1B: out_word = 8'hEB;
		16'hDF1C: out_word = 8'hC9;
		16'hDF1D: out_word = 8'hFF;
		16'hDF1E: out_word = 8'h11;
		16'hDF1F: out_word = 8'hEA;
		16'hDF20: out_word = 8'h6B;
		16'hDF21: out_word = 8'h26;
		16'hDF22: out_word = 8'h0A;
		16'hDF23: out_word = 8'h06;
		16'hDF24: out_word = 8'h08;
		16'hDF25: out_word = 8'hEB;
		16'hDF26: out_word = 8'hC5;
		16'hDF27: out_word = 8'h5E;
		16'hDF28: out_word = 8'h23;
		16'hDF29: out_word = 8'h4F;
		16'hDF2A: out_word = 8'h91;
		16'hDF2B: out_word = 8'h24;
		16'hDF2C: out_word = 8'h10;
		16'hDF2D: out_word = 8'hF6;
		16'hDF2E: out_word = 8'hC9;
		16'hDF2F: out_word = 8'hFF;
		16'hDF30: out_word = 8'h3A;
		16'hDF31: out_word = 8'h55;
		16'hDF32: out_word = 8'h6C;
		16'hDF33: out_word = 8'hE6;
		16'hDF34: out_word = 8'h04;
		16'hDF35: out_word = 8'hC8;
		16'hDF36: out_word = 8'h26;
		16'hDF37: out_word = 8'h0C;
		16'hDF38: out_word = 8'h40;
		16'hDF39: out_word = 8'h94;
		16'hDF3A: out_word = 8'h26;
		16'hDF3B: out_word = 8'h10;
		16'hDF3C: out_word = 8'hF8;
		16'hDF3D: out_word = 8'h11;
		16'hDF3E: out_word = 8'h99;
		16'hDF3F: out_word = 8'hF8;
		16'hDF40: out_word = 8'hFE;
		16'hDF41: out_word = 8'h55;
		16'hDF42: out_word = 8'h7E;
		16'hDF43: out_word = 8'hE6;
		16'hDF44: out_word = 8'hD9;
		16'hDF45: out_word = 8'h01;
		16'hDF46: out_word = 8'h22;
		16'hDF47: out_word = 8'hD6;
		16'hDF48: out_word = 8'h04;
		16'hDF49: out_word = 8'h82;
		16'hDF4A: out_word = 8'hF3;
		16'hDF4B: out_word = 8'hFF;
		16'hDF4C: out_word = 8'h24;
		16'hDF4D: out_word = 8'h83;
		16'hDF4E: out_word = 8'h0A;
		16'hDF4F: out_word = 8'hEE;
		16'hDF50: out_word = 8'h1A;
		16'hDF51: out_word = 8'h02;
		16'hDF52: out_word = 8'h03;
		16'hDF53: out_word = 8'h8A;
		16'hDF54: out_word = 8'h26;
		16'hDF55: out_word = 8'hCA;
		16'hDF56: out_word = 8'h5A;
		16'hDF57: out_word = 8'hF3;
		16'hDF58: out_word = 8'h00;
		16'hDF59: out_word = 8'h33;
		16'hDF5A: out_word = 8'hF3;
		16'hDF5B: out_word = 8'h01;
		16'hDF5C: out_word = 8'h2D;
		16'hDF5D: out_word = 8'hDB;
		16'hDF5E: out_word = 8'h07;
		16'hDF5F: out_word = 8'h68;
		16'hDF60: out_word = 8'hF5;
		16'hDF61: out_word = 8'h36;
		16'hDF62: out_word = 8'hEC;
		16'hDF63: out_word = 8'h08;
		16'hDF64: out_word = 8'hCB;
		16'hDF65: out_word = 8'hF7;
		16'hDF66: out_word = 8'h09;
		16'hDF67: out_word = 8'h47;
		16'hDF68: out_word = 8'hF7;
		16'hDF69: out_word = 8'h21;
		16'hDF6A: out_word = 8'h1D;
		16'hDF6B: out_word = 8'h6B;
		16'hDF6C: out_word = 8'h58;
		16'hDF6D: out_word = 8'h64;
		16'hDF6E: out_word = 8'hEB;
		16'hDF6F: out_word = 8'hD9;
		16'hDF70: out_word = 8'hC9;
		16'hDF71: out_word = 8'hE5;
		16'hDF72: out_word = 8'hD8;
		16'hDF73: out_word = 8'h15;
		16'hDF74: out_word = 8'h11;
		16'hDF75: out_word = 8'h0A;
		16'hDF76: out_word = 8'hBD;
		16'hDF77: out_word = 8'hAF;
		16'hDF78: out_word = 8'h3D;
		16'hDF79: out_word = 8'h3C;
		16'hDF7A: out_word = 8'hD6;
		16'hDF7B: out_word = 8'hB1;
		16'hDF7C: out_word = 8'hC4;
		16'hDF7D: out_word = 8'h19;
		16'hDF7E: out_word = 8'hC6;
		16'hDF7F: out_word = 8'hCF;
		16'hDF80: out_word = 8'h57;
		16'hDF81: out_word = 8'h7D;
		16'hDF82: out_word = 8'hFC;
		16'hDF83: out_word = 8'hE1;
		16'hDF84: out_word = 8'h72;
		16'hDF85: out_word = 8'h23;
		16'hDF86: out_word = 8'h8D;
		16'hDF87: out_word = 8'h77;
		16'hDF88: out_word = 8'hC9;
		16'hDF89: out_word = 8'h59;
		16'hDF8A: out_word = 8'hB7;
		16'hDF8B: out_word = 8'h5B;
		16'hDF8C: out_word = 8'hD3;
		16'hDF8D: out_word = 8'h6E;
		16'hDF8E: out_word = 8'hE7;
		16'hDF8F: out_word = 8'h30;
		16'hDF90: out_word = 8'hA7;
		16'hDF91: out_word = 8'h3E;
		16'hDF92: out_word = 8'h27;
		16'hDF93: out_word = 8'h85;
		16'hDF94: out_word = 8'hFB;
		16'hDF95: out_word = 8'hC9;
		16'hDF96: out_word = 8'hF3;
		16'hDF97: out_word = 8'hFF;
		16'hDF98: out_word = 8'hDD;
		16'hDF99: out_word = 8'h21;
		16'hDF9A: out_word = 8'hC1;
		16'hDF9B: out_word = 8'h2F;
		16'hDF9C: out_word = 8'hCD;
		16'hDF9D: out_word = 8'h26;
		16'hDF9E: out_word = 8'h86;
		16'hDF9F: out_word = 8'h3E;
		16'hDFA0: out_word = 8'hE7;
		16'hDFA1: out_word = 8'h08;
		16'hDFA2: out_word = 8'h0E;
		16'hDFA3: out_word = 8'h1F;
		16'hDFA4: out_word = 8'hF5;
		16'hDFA5: out_word = 8'h53;
		16'hDFA6: out_word = 8'h2A;
		16'hDFA7: out_word = 8'h4D;
		16'hDFA8: out_word = 8'hF5;
		16'hDFA9: out_word = 8'h06;
		16'hDFAA: out_word = 8'h00;
		16'hDFAB: out_word = 8'h4F;
		16'hDFAC: out_word = 8'hB5;
		16'hDFAD: out_word = 8'hD8;
		16'hDFAE: out_word = 8'h5C;
		16'hDFAF: out_word = 8'hFF;
		16'hDFB0: out_word = 8'hCD;
		16'hDFB1: out_word = 8'h77;
		16'hDFB2: out_word = 8'h83;
		16'hDFB3: out_word = 8'hF5;
		16'hDFB4: out_word = 8'h3E;
		16'hDFB5: out_word = 8'hC9;
		16'hDFB6: out_word = 8'h32;
		16'hDFB7: out_word = 8'hC2;
		16'hDFB8: out_word = 8'hCC;
		16'hDFB9: out_word = 8'h5C;
		16'hDFBA: out_word = 8'hAF;
		16'hDFBB: out_word = 8'hE8;
		16'hDFBC: out_word = 8'hF3;
		16'hDFBD: out_word = 8'hBA;
		16'hDFBE: out_word = 8'h01;
		16'hDFBF: out_word = 8'h77;
		16'hDFC0: out_word = 8'hCF;
		16'hDFC1: out_word = 8'hEB;
		16'hDFC2: out_word = 8'h1A;
		16'hDFC3: out_word = 8'hF9;
		16'hDFC4: out_word = 8'hBF;
		16'hDFC5: out_word = 8'hCF;
		16'hDFC6: out_word = 8'hF1;
		16'hDFC7: out_word = 8'hFB;
		16'hDFC8: out_word = 8'hC9;
		16'hDFC9: out_word = 8'hED;
		16'hDFCA: out_word = 8'h73;
		16'hDFCB: out_word = 8'h8E;
		16'hDFCC: out_word = 8'hE9;
		16'hDFCD: out_word = 8'h83;
		16'hDFCE: out_word = 8'h3E;
		16'hDFCF: out_word = 8'hC3;
		16'hDFD0: out_word = 8'hDE;
		16'hDFD1: out_word = 8'h21;
		16'hDFD2: out_word = 8'h81;
		16'hDFD3: out_word = 8'h8D;
		16'hDFD4: out_word = 8'h22;
		16'hDFD5: out_word = 8'h00;
		16'hDFD6: out_word = 8'h25;
		16'hDFD7: out_word = 8'h3A;
		16'hDFD8: out_word = 8'h57;
		16'hDFD9: out_word = 8'h20;
		16'hDFDA: out_word = 8'h9D;
		16'hDFDB: out_word = 8'hA8;
		16'hDFDC: out_word = 8'h31;
		16'hDFDD: out_word = 8'h5C;
		16'hDFDE: out_word = 8'h18;
		16'hDFDF: out_word = 8'hFF;
		16'hDFE0: out_word = 8'h15;
		16'hDFE1: out_word = 8'h51;
		16'hDFE2: out_word = 8'h6C;
		16'hDFE3: out_word = 8'hA7;
		16'hDFE4: out_word = 8'hC8;
		16'hDFE5: out_word = 8'hDD;
		16'hDFE6: out_word = 8'hE5;
		16'hDFE7: out_word = 8'hCD;
		16'hDFE8: out_word = 8'hC3;
		16'hDFE9: out_word = 8'h3B;
		16'hDFEA: out_word = 8'h83;
		16'hDFEB: out_word = 8'hFC;
		16'hDFEC: out_word = 8'hE1;
		16'hDFED: out_word = 8'h21;
		16'hDFEE: out_word = 8'h52;
		16'hDFEF: out_word = 8'h6C;
		16'hDFF0: out_word = 8'hBE;
		16'hDFF1: out_word = 8'hC8;
		16'hDFF2: out_word = 8'h25;
		16'hDFF3: out_word = 8'h36;
		16'hDFF4: out_word = 8'h66;
		16'hDFF5: out_word = 8'h8D;
		16'hDFF6: out_word = 8'hD4;
		16'hDFF7: out_word = 8'hB7;
		16'hDFF8: out_word = 8'h85;
		16'hDFF9: out_word = 8'h1D;
		16'hDFFA: out_word = 8'hD4;
		16'hDFFB: out_word = 8'hEB;
		16'hDFFC: out_word = 8'h05;
		16'hDFFD: out_word = 8'h9E;
		16'hDFFE: out_word = 8'hA5;
		16'hDFFF: out_word = 8'hCA;
		16'hE000: out_word = 8'h08;
		16'hE001: out_word = 8'h13;
		16'hE002: out_word = 8'h01;
		16'hE003: out_word = 8'h05;
		16'hE004: out_word = 8'h19;
		16'hE005: out_word = 8'h53;
		16'hE006: out_word = 8'h84;
		16'hE007: out_word = 8'h3A;
		16'hE008: out_word = 8'hE7;
		16'hE009: out_word = 8'hF0;
		16'hE00A: out_word = 8'hC0;
		16'hE00B: out_word = 8'hFE;
		16'hE00C: out_word = 8'h10;
		16'hE00D: out_word = 8'hC2;
		16'hE00E: out_word = 8'hEF;
		16'hE00F: out_word = 8'h75;
		16'hE010: out_word = 8'h92;
		16'hE011: out_word = 8'hB6;
		16'hE012: out_word = 8'h5E;
		16'hE013: out_word = 8'hEC;
		16'hE014: out_word = 8'h09;
		16'hE015: out_word = 8'hEC;
		16'hE016: out_word = 8'hA5;
		16'hE017: out_word = 8'hC8;
		16'hE018: out_word = 8'hEC;
		16'hE019: out_word = 8'hF0;
		16'hE01A: out_word = 8'h4C;
		16'hE01B: out_word = 8'h08;
		16'hE01C: out_word = 8'hA7;
		16'hE01D: out_word = 8'hEB;
		16'hE01E: out_word = 8'h41;
		16'hE01F: out_word = 8'h3A;
		16'hE020: out_word = 8'hE4;
		16'hE021: out_word = 8'hC8;
		16'hE022: out_word = 8'hC2;
		16'hE023: out_word = 8'h47;
		16'hE024: out_word = 8'h0E;
		16'hE025: out_word = 8'h99;
		16'hE026: out_word = 8'hD9;
		16'hE027: out_word = 8'hAA;
		16'hE028: out_word = 8'hD1;
		16'hE029: out_word = 8'hFC;
		16'hE02A: out_word = 8'hFD;
		16'hE02B: out_word = 8'h7E;
		16'hE02C: out_word = 8'h08;
		16'hE02D: out_word = 8'hFE;
		16'hE02E: out_word = 8'h42;
		16'hE02F: out_word = 8'h20;
		16'hE030: out_word = 8'h2C;
		16'hE031: out_word = 8'h7B;
		16'hE032: out_word = 8'h94;
		16'hE033: out_word = 8'h3D;
		16'hE034: out_word = 8'h28;
		16'hE035: out_word = 8'hA5;
		16'hE036: out_word = 8'h26;
		16'hE037: out_word = 8'hEE;
		16'hE038: out_word = 8'hE1;
		16'hE039: out_word = 8'h8F;
		16'hE03A: out_word = 8'h67;
		16'hE03B: out_word = 8'h7E;
		16'hE03C: out_word = 8'hD9;
		16'hE03D: out_word = 8'h0C;
		16'hE03E: out_word = 8'h58;
		16'hE03F: out_word = 8'hE7;
		16'hE040: out_word = 8'h53;
		16'hE041: out_word = 8'h8E;
		16'hE042: out_word = 8'hC0;
		16'hE043: out_word = 8'h92;
		16'hE044: out_word = 8'h68;
		16'hE045: out_word = 8'hE0;
		16'hE046: out_word = 8'h36;
		16'hE047: out_word = 8'h0F;
		16'hE048: out_word = 8'h00;
		16'hE049: out_word = 8'h60;
		16'hE04A: out_word = 8'h71;
		16'hE04B: out_word = 8'h10;
		16'hE04C: out_word = 8'hE6;
		16'hE04D: out_word = 8'h70;
		16'hE04E: out_word = 8'h11;
		16'hE04F: out_word = 8'hF6;
		16'hE050: out_word = 8'h12;
		16'hE051: out_word = 8'h44;
		16'hE052: out_word = 8'hF6;
		16'hE053: out_word = 8'h89;
		16'hE054: out_word = 8'h13;
		16'hE055: out_word = 8'h78;
		16'hE056: out_word = 8'hF5;
		16'hE057: out_word = 8'hB1;
		16'hE058: out_word = 8'hCA;
		16'hE059: out_word = 8'h06;
		16'hE05A: out_word = 8'h85;
		16'hE05B: out_word = 8'hCF;
		16'hE05C: out_word = 8'h93;
		16'hE05D: out_word = 8'h96;
		16'hE05E: out_word = 8'h78;
		16'hE05F: out_word = 8'hA7;
		16'hE060: out_word = 8'h79;
		16'hE061: out_word = 8'hFD;
		16'hE062: out_word = 8'h20;
		16'hE063: out_word = 8'h0A;
		16'hE064: out_word = 8'hFE;
		16'hE065: out_word = 8'h17;
		16'hE066: out_word = 8'h38;
		16'hE067: out_word = 8'h06;
		16'hE068: out_word = 8'h3F;
		16'hE069: out_word = 8'hF3;
		16'hE06A: out_word = 8'hD6;
		16'hE06B: out_word = 8'h3E;
		16'hE06C: out_word = 8'h16;
		16'hE06D: out_word = 8'h32;
		16'hE06E: out_word = 8'hCF;
		16'hE06F: out_word = 8'h84;
		16'hE070: out_word = 8'hF1;
		16'hE071: out_word = 8'hC6;
		16'hE072: out_word = 8'h02;
		16'hE073: out_word = 8'hDD;
		16'hE074: out_word = 8'h77;
		16'hE075: out_word = 8'h4E;
		16'hE076: out_word = 8'hDC;
		16'hE077: out_word = 8'h03;
		16'hE078: out_word = 8'h0C;
		16'hE079: out_word = 8'hFE;
		16'hE07A: out_word = 8'hFD;
		16'hE07B: out_word = 8'h55;
		16'hE07C: out_word = 8'h28;
		16'hE07D: out_word = 8'h14;
		16'hE07E: out_word = 8'hDD;
		16'hE07F: out_word = 8'h34;
		16'hE080: out_word = 8'h03;
		16'hE081: out_word = 8'h7A;
		16'hE082: out_word = 8'h2F;
		16'hE083: out_word = 8'hF5;
		16'hE084: out_word = 8'h44;
		16'hE085: out_word = 8'hEE;
		16'hE086: out_word = 8'hA9;
		16'hE087: out_word = 8'h18;
		16'hE088: out_word = 8'hD0;
		16'hE089: out_word = 8'h46;
		16'hE08A: out_word = 8'hF1;
		16'hE08B: out_word = 8'hE3;
		16'hE08C: out_word = 8'h0A;
		16'hE08D: out_word = 8'h03;
		16'hE08E: out_word = 8'h2F;
		16'hE08F: out_word = 8'hF7;
		16'hE090: out_word = 8'h29;
		16'hE091: out_word = 8'h06;
		16'hE092: out_word = 8'h35;
		16'hE093: out_word = 8'hB9;
		16'hE094: out_word = 8'hEF;
		16'hE095: out_word = 8'hB9;
		16'hE096: out_word = 8'h5E;
		16'hE097: out_word = 8'h0F;
		16'hE098: out_word = 8'hAF;
		16'hE099: out_word = 8'hEA;
		16'hE09A: out_word = 8'h57;
		16'hE09B: out_word = 8'hED;
		16'hE09C: out_word = 8'h52;
		16'hE09D: out_word = 8'h37;
		16'hE09E: out_word = 8'hA8;
		16'hE09F: out_word = 8'h29;
		16'hE0A0: out_word = 8'h7F;
		16'hE0A1: out_word = 8'h10;
		16'hE0A2: out_word = 8'h08;
		16'hE0A3: out_word = 8'h20;
		16'hE0A4: out_word = 8'hBB;
		16'hE0A5: out_word = 8'h26;
		16'hE0A6: out_word = 8'h4A;
		16'hE0A7: out_word = 8'h5F;
		16'hE0A8: out_word = 8'hD1;
		16'hE0A9: out_word = 8'h34;
		16'hE0AA: out_word = 8'h0D;
		16'hE0AB: out_word = 8'hDA;
		16'hE0AC: out_word = 8'h6A;
		16'hE0AD: out_word = 8'h3E;
		16'hE0AE: out_word = 8'h14;
		16'hE0AF: out_word = 8'h3F;
		16'hE0B0: out_word = 8'h1C;
		16'hE0B1: out_word = 8'h06;
		16'hE0B2: out_word = 8'h08;
		16'hE0B3: out_word = 8'hB5;
		16'hE0B4: out_word = 8'hD5;
		16'hE0B5: out_word = 8'hEA;
		16'hE0B6: out_word = 8'h1B;
		16'hE0B7: out_word = 8'h7F;
		16'hE0B8: out_word = 8'h00;
		16'hE0B9: out_word = 8'h19;
		16'hE0BA: out_word = 8'hD1;
		16'hE0BB: out_word = 8'h1C;
		16'hE0BC: out_word = 8'h0D;
		16'hE0BD: out_word = 8'h20;
		16'hE0BE: out_word = 8'hED;
		16'hE0BF: out_word = 8'hC9;
		16'hE0C0: out_word = 8'h05;
		16'hE0C1: out_word = 8'hB8;
		16'hE0C2: out_word = 8'hE2;
		16'hE0C3: out_word = 8'hD7;
		16'hE0C4: out_word = 8'h1C;
		16'hE0C5: out_word = 8'hC5;
		16'hE0C6: out_word = 8'h86;
		16'hE0C7: out_word = 8'h89;
		16'hE0C8: out_word = 8'hB2;
		16'hE0C9: out_word = 8'hE5;
		16'hE0CA: out_word = 8'h7B;
		16'hE0CB: out_word = 8'h07;
		16'hE0CC: out_word = 8'hD1;
		16'hE0CD: out_word = 8'hB3;
		16'hE0CE: out_word = 8'hD5;
		16'hE0CF: out_word = 8'h7A;
		16'hE0D0: out_word = 8'h05;
		16'hE0D1: out_word = 8'hBA;
		16'hE0D2: out_word = 8'h06;
		16'hE0D3: out_word = 8'hDF;
		16'hE0D4: out_word = 8'h9D;
		16'hE0D5: out_word = 8'hD7;
		16'hE0D6: out_word = 8'hD1;
		16'hE0D7: out_word = 8'hE1;
		16'hE0D8: out_word = 8'hC1;
		16'hE0D9: out_word = 8'h29;
		16'hE0DA: out_word = 8'hBE;
		16'hE0DB: out_word = 8'hCB;
		16'hE0DC: out_word = 8'h22;
		16'hE0DD: out_word = 8'h1E;
		16'hE0DE: out_word = 8'hB4;
		16'hE0DF: out_word = 8'h69;
		16'hE0E0: out_word = 8'h94;
		16'hE0E1: out_word = 8'h2F;
		16'hE0E2: out_word = 8'hF3;
		16'hE0E3: out_word = 8'h1D;
		16'hE0E4: out_word = 8'h59;
		16'hE0E5: out_word = 8'h63;
		16'hE0E6: out_word = 8'hA1;
		16'hE0E7: out_word = 8'h72;
		16'hE0E8: out_word = 8'hC7;
		16'hE0E9: out_word = 8'h79;
		16'hE0EA: out_word = 8'h00;
		16'hE0EB: out_word = 8'h80;
		16'hE0EC: out_word = 8'hF7;
		16'hE0ED: out_word = 8'h73;
		16'hE0EE: out_word = 8'h6C;
		16'hE0EF: out_word = 8'h01;
		16'hE0F0: out_word = 8'h08;
		16'hE0F1: out_word = 8'h47;
		16'hE0F2: out_word = 8'h24;
		16'hE0F3: out_word = 8'hAF;
		16'hE0F4: out_word = 8'h3E;
		16'hE0F5: out_word = 8'hC7;
		16'hE0F6: out_word = 8'h11;
		16'hE0F7: out_word = 8'hFF;
		16'hE0F8: out_word = 8'hFF;
		16'hE0F9: out_word = 8'h0E;
		16'hE0FA: out_word = 8'hA8;
		16'hE0FB: out_word = 8'hED;
		16'hE0FC: out_word = 8'hB8;
		16'hE0FD: out_word = 8'h21;
		16'hE0FE: out_word = 8'h56;
		16'hE0FF: out_word = 8'h6C;
		16'hE100: out_word = 8'h11;
		16'hE101: out_word = 8'hF4;
		16'hE102: out_word = 8'h3B;
		16'hE103: out_word = 8'h5D;
		16'hE104: out_word = 8'h01;
		16'hE105: out_word = 8'h28;
		16'hE106: out_word = 8'hEB;
		16'hE107: out_word = 8'h51;
		16'hE108: out_word = 8'hEC;
		16'hE109: out_word = 8'hF1;
		16'hE10A: out_word = 8'hFD;
		16'hE10B: out_word = 8'h21;
		16'hE10C: out_word = 8'h3A;
		16'hE10D: out_word = 8'h5C;
		16'hE10E: out_word = 8'h39;
		16'hE10F: out_word = 8'h36;
		16'hE110: out_word = 8'h00;
		16'hE111: out_word = 8'hFF;
		16'hE112: out_word = 8'h06;
		16'hE113: out_word = 8'hD3;
		16'hE114: out_word = 8'h01;
		16'hE115: out_word = 8'hFE;
		16'hE116: out_word = 8'hFC;
		16'hE117: out_word = 8'hA6;
		16'hE118: out_word = 8'h21;
		16'hE119: out_word = 8'hEF;
		16'hE11A: out_word = 8'h58;
		16'hE11B: out_word = 8'h27;
		16'hE11C: out_word = 8'hD9;
		16'hE11D: out_word = 8'hFF;
		16'hE11E: out_word = 8'h03;
		16'hE11F: out_word = 8'h21;
		16'hE120: out_word = 8'h01;
		16'hE121: out_word = 8'h00;
		16'hE122: out_word = 8'hC2;
		16'hE123: out_word = 8'h22;
		16'hE124: out_word = 8'h42;
		16'hE125: out_word = 8'hE2;
		16'hE126: out_word = 8'hAF;
		16'hE127: out_word = 8'h32;
		16'hE128: out_word = 8'h44;
		16'hE129: out_word = 8'h7E;
		16'hE12A: out_word = 8'h01;
		16'hE12B: out_word = 8'hFF;
		16'hE12C: out_word = 8'h5F;
		16'hE12D: out_word = 8'hCD;
		16'hE12E: out_word = 8'hB7;
		16'hE12F: out_word = 8'h1E;
		16'hE130: out_word = 8'hE8;
		16'hE131: out_word = 8'h7F;
		16'hE132: out_word = 8'hE7;
		16'hE133: out_word = 8'hFB;
		16'hE134: out_word = 8'hC3;
		16'hE135: out_word = 8'h7D;
		16'hE136: out_word = 8'h1B;
		16'hE137: out_word = 8'h3A;
		16'hE138: out_word = 8'hE9;
		16'hE139: out_word = 8'h6A;
		16'hE13A: out_word = 8'hFE;
		16'hE13B: out_word = 8'h3C;
		16'hE13C: out_word = 8'hD6;
		16'hE13D: out_word = 8'h10;
		16'hE13E: out_word = 8'hFE;
		16'hE13F: out_word = 8'h35;
		16'hE140: out_word = 8'h38;
		16'hE141: out_word = 8'h07;
		16'hE142: out_word = 8'h17;
		16'hE143: out_word = 8'h04;
		16'hE144: out_word = 8'h18;
		16'hE145: out_word = 8'h03;
		16'hE146: out_word = 8'h7C;
		16'hE147: out_word = 8'hBF;
		16'hE148: out_word = 8'h9F;
		16'hE149: out_word = 8'h21;
		16'hE14A: out_word = 8'hD8;
		16'hE14B: out_word = 8'h60;
		16'hE14C: out_word = 8'hE5;
		16'hE14D: out_word = 8'h32;
		16'hE14E: out_word = 8'h50;
		16'hE14F: out_word = 8'hDA;
		16'hE150: out_word = 8'h6C;
		16'hE151: out_word = 8'h6F;
		16'hE152: out_word = 8'hFA;
		16'hE153: out_word = 8'h19;
		16'hE154: out_word = 8'h10;
		16'hE155: out_word = 8'hEE;
		16'hE156: out_word = 8'hEE;
		16'hE157: out_word = 8'h9B;
		16'hE158: out_word = 8'h1F;
		16'hE159: out_word = 8'h63;
		16'hE15A: out_word = 8'hE6;
		16'hE15B: out_word = 8'hE7;
		16'hE15C: out_word = 8'h60;
		16'hE15D: out_word = 8'h62;
		16'hE15E: out_word = 8'hB8;
		16'hE15F: out_word = 8'hE7;
		16'hE160: out_word = 8'hE7;
		16'hE161: out_word = 8'hE9;
		16'hE162: out_word = 8'h02;
		16'hE163: out_word = 8'h28;
		16'hE164: out_word = 8'h08;
		16'hE165: out_word = 8'hFF;
		16'hE166: out_word = 8'h3E;
		16'hE167: out_word = 8'hFA;
		16'hE168: out_word = 8'hDB;
		16'hE169: out_word = 8'hDF;
		16'hE16A: out_word = 8'h1F;
		16'hE16B: out_word = 8'hD2;
		16'hE16C: out_word = 8'hF0;
		16'hE16D: out_word = 8'h75;
		16'hE16E: out_word = 8'hE3;
		16'hE16F: out_word = 8'hF1;
		16'hE170: out_word = 8'hE3;
		16'hE171: out_word = 8'hC9;
		16'hE172: out_word = 8'h6B;
		16'hE173: out_word = 8'hF5;
		16'hE174: out_word = 8'h7C;
		16'hE175: out_word = 8'h18;
		16'hE176: out_word = 8'hE3;
		16'hE177: out_word = 8'hE7;
		16'hE178: out_word = 8'h7D;
		16'hE179: out_word = 8'h70;
		16'hE17A: out_word = 8'h6B;
		16'hE17B: out_word = 8'hF7;
		16'hE17C: out_word = 8'hE2;
		16'hE17D: out_word = 8'hE1;
		16'hE17E: out_word = 8'h2B;
		16'hE17F: out_word = 8'hFF;
		16'hE180: out_word = 8'hFB;
		16'hE181: out_word = 8'hDF;
		16'hE182: out_word = 8'hDB;
		16'hE183: out_word = 8'h21;
		16'hE184: out_word = 8'hF4;
		16'hE185: out_word = 8'h5C;
		16'hE186: out_word = 8'h7E;
		16'hE187: out_word = 8'h3C;
		16'hE188: out_word = 8'h03;
		16'hE189: out_word = 8'h49;
		16'hE18A: out_word = 8'h86;
		16'hE18B: out_word = 8'hF1;
		16'hE18C: out_word = 8'h32;
		16'hE18D: out_word = 8'h77;
		16'hE18E: out_word = 8'h65;
		16'hE18F: out_word = 8'h7A;
		16'hE190: out_word = 8'h22;
		16'hE191: out_word = 8'h76;
		16'hE192: out_word = 8'h7F;
		16'hE193: out_word = 8'h23;
		16'hE194: out_word = 8'h7E;
		16'hE195: out_word = 8'hCB;
		16'hE196: out_word = 8'h3F;
		16'hE197: out_word = 8'h5F;
		16'hE198: out_word = 8'hCE;
		16'hE199: out_word = 8'h30;
		16'hE19A: out_word = 8'hFB;
		16'hE19B: out_word = 8'h93;
		16'hE19C: out_word = 8'h32;
		16'hE19D: out_word = 8'h79;
		16'hE19E: out_word = 8'h65;
		16'hE19F: out_word = 8'h7B;
		16'hE1A0: out_word = 8'h94;
		16'hE1A1: out_word = 8'hEA;
		16'hE1A2: out_word = 8'h74;
		16'hE1A3: out_word = 8'hEA;
		16'hE1A4: out_word = 8'h88;
		16'hE1A5: out_word = 8'h73;
		16'hE1A6: out_word = 8'h6D;
		16'hE1A7: out_word = 8'h15;
		16'hE1A8: out_word = 8'h40;
		16'hE1A9: out_word = 8'h63;
		16'hE1AA: out_word = 8'h44;
		16'hE1AB: out_word = 8'h0E;
		16'hE1AC: out_word = 8'hDA;
		16'hE1AD: out_word = 8'hFF;
		16'hE1AE: out_word = 8'hAF;
		16'hE1AF: out_word = 8'hF9;
		16'hE1B0: out_word = 8'h49;
		16'hE1B1: out_word = 8'h4B;
		16'hE1B2: out_word = 8'h0B;
		16'hE1B3: out_word = 8'hF6;
		16'hE1B4: out_word = 8'h3C;
		16'hE1B5: out_word = 8'h77;
		16'hE1B6: out_word = 8'hB7;
		16'hE1B7: out_word = 8'h36;
		16'hE1B8: out_word = 8'h68;
		16'hE1B9: out_word = 8'h0E;
		16'hE1BA: out_word = 8'h7B;
		16'hE1BB: out_word = 8'h59;
		16'hE1BC: out_word = 8'h21;
		16'hE1BD: out_word = 8'h9D;
		16'hE1BE: out_word = 8'hCB;
		16'hE1BF: out_word = 8'h65;
		16'hE1C0: out_word = 8'h22;
		16'hE1C1: out_word = 8'h55;
		16'hE1C2: out_word = 8'h27;
		16'hE1C3: out_word = 8'hDD;
		16'hE1C4: out_word = 8'h8D;
		16'hE1C5: out_word = 8'hC9;
		16'hE1C6: out_word = 8'hDD;
		16'hE1C7: out_word = 8'hE5;
		16'hE1C8: out_word = 8'h40;
		16'hE1C9: out_word = 8'h03;
		16'hE1CA: out_word = 8'hFE;
		16'hE1CB: out_word = 8'hB2;
		16'hE1CC: out_word = 8'h32;
		16'hE1CD: out_word = 8'h42;
		16'hE1CE: out_word = 8'h86;
		16'hE1CF: out_word = 8'h17;
		16'hE1D0: out_word = 8'h0E;
		16'hE1D1: out_word = 8'h02;
		16'hE1D2: out_word = 8'hBC;
		16'hE1D3: out_word = 8'hA1;
		16'hE1D4: out_word = 8'hFF;
		16'hE1D5: out_word = 8'h66;
		16'hE1D6: out_word = 8'h1A;
		16'hE1D7: out_word = 8'h21;
		16'hE1D8: out_word = 8'h0F;
		16'hE1D9: out_word = 8'hD9;
		16'hE1DA: out_word = 8'hE6;
		16'hE1DB: out_word = 8'h15;
		16'hE1DC: out_word = 8'h1E;
		16'hE1DD: out_word = 8'h53;
		16'hE1DE: out_word = 8'hB6;
		16'hE1DF: out_word = 8'hFD;
		16'hE1E0: out_word = 8'h1F;
		16'hE1E1: out_word = 8'h87;
		16'hE1E2: out_word = 8'h18;
		16'hE1E3: out_word = 8'h16;
		16'hE1E4: out_word = 8'hFF;
		16'hE1E5: out_word = 8'h2F;
		16'hE1E6: out_word = 8'h14;
		16'hE1E7: out_word = 8'hD6;
		16'hE1E8: out_word = 8'h0A;
		16'hE1E9: out_word = 8'h30;
		16'hE1EA: out_word = 8'hFB;
		16'hE1EB: out_word = 8'hC6;
		16'hE1EC: out_word = 8'h3A;
		16'hE1ED: out_word = 8'hEA;
		16'hE1EE: out_word = 8'hC9;
		16'hE1EF: out_word = 8'h3E;
		16'hE1F0: out_word = 8'h52;
		16'hE1F1: out_word = 8'h1F;
		16'hE1F2: out_word = 8'hF1;
		16'hE1F3: out_word = 8'h49;
		16'hE1F4: out_word = 8'h21;
		16'hE1F5: out_word = 8'h7E;
		16'hE1F6: out_word = 8'h3F;
		16'hE1F7: out_word = 8'hE3;
		16'hE1F8: out_word = 8'hA7;
		16'hE1F9: out_word = 8'hF3;
		16'hE1FA: out_word = 8'hCA;
		16'hE1FB: out_word = 8'hF5;
		16'hE1FC: out_word = 8'h87;
		16'hE1FD: out_word = 8'h6F;
		16'hE1FE: out_word = 8'hF7;
		16'hE1FF: out_word = 8'h5F;
		16'hE200: out_word = 8'h26;
		16'hE201: out_word = 8'h00;
		16'hE202: out_word = 8'h54;
		16'hE203: out_word = 8'h7C;
		16'hE204: out_word = 8'hB6;
		16'hE205: out_word = 8'hF0;
		16'hE206: out_word = 8'hFD;
		16'hE207: out_word = 8'h11;
		16'hE208: out_word = 8'h90;
		16'hE209: out_word = 8'h6C;
		16'hE20A: out_word = 8'h84;
		16'hE20B: out_word = 8'hF5;
		16'hE20C: out_word = 8'h5C;
		16'hE20D: out_word = 8'h50;
		16'hE20E: out_word = 8'h0E;
		16'hE20F: out_word = 8'h03;
		16'hE210: out_word = 8'hFE;
		16'hE211: out_word = 8'h7E;
		16'hE212: out_word = 8'h12;
		16'hE213: out_word = 8'h23;
		16'hE214: out_word = 8'h1C;
		16'hE215: out_word = 8'hD5;
		16'hE216: out_word = 8'hFC;
		16'hE217: out_word = 8'h1D;
		16'hE218: out_word = 8'h1F;
		16'hE219: out_word = 8'h14;
		16'hE21A: out_word = 8'h10;
		16'hE21B: out_word = 8'hBA;
		16'hE21C: out_word = 8'hF0;
		16'hE21D: out_word = 8'h8E;
		16'hE21E: out_word = 8'hF8;
		16'hE21F: out_word = 8'hA1;
		16'hE220: out_word = 8'hFA;
		16'hE221: out_word = 8'h2A;
		16'hE222: out_word = 8'hE3;
		16'hE223: out_word = 8'hE3;
		16'hE224: out_word = 8'h21;
		16'hE225: out_word = 8'h47;
		16'hE226: out_word = 8'hF1;
		16'hE227: out_word = 8'h22;
		16'hE228: out_word = 8'h5C;
		16'hE229: out_word = 8'h5A;
		16'hE22A: out_word = 8'h66;
		16'hE22B: out_word = 8'h5D;
		16'hE22C: out_word = 8'hFD;
		16'hE22D: out_word = 8'h7C;
		16'hE22E: out_word = 8'h66;
		16'hE22F: out_word = 8'hFD;
		16'hE230: out_word = 8'h7D;
		16'hE231: out_word = 8'hFD;
		16'hE232: out_word = 8'h9C;
		16'hE233: out_word = 8'h61;
		16'hE234: out_word = 8'hFD;
		16'hE235: out_word = 8'h9D;
		16'hE236: out_word = 8'h75;
		16'hE237: out_word = 8'hF1;
		16'hE238: out_word = 8'hC9;
		16'hE239: out_word = 8'hF5;
		16'hE23A: out_word = 8'hEF;
		16'hE23B: out_word = 8'hA4;
		16'hE23C: out_word = 8'h5E;
		16'hE23D: out_word = 8'h28;
		16'hE23E: out_word = 8'h2A;
		16'hE23F: out_word = 8'h3A;
		16'hE240: out_word = 8'hF3;
		16'hE241: out_word = 8'h8E;
		16'hE242: out_word = 8'h6C;
		16'hE243: out_word = 8'h3C;
		16'hE244: out_word = 8'h32;
		16'hE245: out_word = 8'hFC;
		16'hE246: out_word = 8'hFE;
		16'hE247: out_word = 8'hF4;
		16'hE248: out_word = 8'h0C;
		16'hE249: out_word = 8'h38;
		16'hE24A: out_word = 8'h35;
		16'hE24B: out_word = 8'hAF;
		16'hE24C: out_word = 8'hF8;
		16'hE24D: out_word = 8'hD0;
		16'hE24E: out_word = 8'h3A;
		16'hE24F: out_word = 8'h8F;
		16'hE250: out_word = 8'hF1;
		16'hE251: out_word = 8'hFF;
		16'hE252: out_word = 8'hFC;
		16'hE253: out_word = 8'hCD;
		16'hE254: out_word = 8'h61;
		16'hE255: out_word = 8'h86;
		16'hE256: out_word = 8'hFE;
		16'hE257: out_word = 8'h09;
		16'hE258: out_word = 8'h38;
		16'hE259: out_word = 8'h23;
		16'hE25A: out_word = 8'hB4;
		16'hE25B: out_word = 8'hAF;
		16'hE25C: out_word = 8'h27;
		16'hE25D: out_word = 8'hF5;
		16'hE25E: out_word = 8'hD6;
		16'hE25F: out_word = 8'h9E;
		16'hE260: out_word = 8'h18;
		16'hE261: out_word = 8'h10;
		16'hE262: out_word = 8'hF9;
		16'hE263: out_word = 8'h2A;
		16'hE264: out_word = 8'h8C;
		16'hE265: out_word = 8'h6C;
		16'hE266: out_word = 8'h23;
		16'hE267: out_word = 8'h22;
		16'hE268: out_word = 8'hFC;
		16'hE269: out_word = 8'hAF;
		16'hE26A: out_word = 8'h7C;
		16'hE26B: out_word = 8'hD2;
		16'hE26C: out_word = 8'hC4;
		16'hE26D: out_word = 8'h0A;
		16'hE26E: out_word = 8'hEE;
		16'hE26F: out_word = 8'hDE;
		16'hE270: out_word = 8'hB0;
		16'hE271: out_word = 8'h16;
		16'hE272: out_word = 8'h85;
		16'hE273: out_word = 8'hF1;
		16'hE274: out_word = 8'hB7;
		16'hE275: out_word = 8'hC2;
		16'hE276: out_word = 8'hE2;
		16'hE277: out_word = 8'hC9;
		16'hE278: out_word = 8'hBB;
		16'hE279: out_word = 8'h9A;
		16'hE27A: out_word = 8'hAF;
		16'hE27B: out_word = 8'hD0;
		16'hE27C: out_word = 8'h67;
		16'hE27D: out_word = 8'h6F;
		16'hE27E: out_word = 8'hEF;
		16'hE27F: out_word = 8'h53;
		16'hE280: out_word = 8'hBB;
		16'hE281: out_word = 8'hC3;
		16'hE282: out_word = 8'h3F;
		16'hE283: out_word = 8'hCD;
		16'hE284: out_word = 8'hE5;
		16'hE285: out_word = 8'h2A;
		16'hE286: out_word = 8'hF0;
		16'hE287: out_word = 8'hCF;
		16'hE288: out_word = 8'hE3;
		16'hE289: out_word = 8'hC5;
		16'hE28A: out_word = 8'hC9;
		16'hE28B: out_word = 8'h08;
		16'hE28C: out_word = 8'hC2;
		16'hE28D: out_word = 8'h7E;
		16'hE28E: out_word = 8'h23;
		16'hE28F: out_word = 8'h98;
		16'hE290: out_word = 8'h87;
		16'hE291: out_word = 8'h11;
		16'hE292: out_word = 8'hFD;
		16'hE293: out_word = 8'hC2;
		16'hE294: out_word = 8'hE0;
		16'hE295: out_word = 8'h21;
		16'hE296: out_word = 8'h2F;
		16'hE297: out_word = 8'h4C;
		16'hE298: out_word = 8'hE3;
		16'hE299: out_word = 8'hFB;
		16'hE29A: out_word = 8'h34;
		16'hE29B: out_word = 8'h3F;
		16'hE29C: out_word = 8'h85;
		16'hE29D: out_word = 8'h6F;
		16'hE29E: out_word = 8'h7C;
		16'hE29F: out_word = 8'hCE;
		16'hE2A0: out_word = 8'hDD;
		16'hE2A1: out_word = 8'h00;
		16'hE2A2: out_word = 8'h67;
		16'hE2A3: out_word = 8'h82;
		16'hE2A4: out_word = 8'h09;
		16'hE2A5: out_word = 8'hE3;
		16'hE2A6: out_word = 8'h71;
		16'hE2A7: out_word = 8'hC5;
		16'hE2A8: out_word = 8'hE1;
		16'hE2A9: out_word = 8'hDD;
		16'hE2AA: out_word = 8'h83;
		16'hE2AB: out_word = 8'hF8;
		16'hE2AC: out_word = 8'h3A;
		16'hE2AD: out_word = 8'h87;
		16'hE2AE: out_word = 8'hEC;
		16'hE2AF: out_word = 8'h88;
		16'hE2B0: out_word = 8'h84;
		16'hE2B1: out_word = 8'h87;
		16'hE2B2: out_word = 8'h95;
		16'hE2B3: out_word = 8'hF2;
		16'hE2B4: out_word = 8'hCF;
		16'hE2B5: out_word = 8'h5D;
		16'hE2B6: out_word = 8'hA1;
		16'hE2B7: out_word = 8'h11;
		16'hE2B8: out_word = 8'h41;
		16'hE2B9: out_word = 8'h5C;
		16'hE2BA: out_word = 8'hF0;
		16'hE2BB: out_word = 8'h5D;
		16'hE2BC: out_word = 8'hE9;
		16'hE2BD: out_word = 8'hA7;
		16'hE2BE: out_word = 8'h3E;
		16'hE2BF: out_word = 8'h06;
		16'hE2C0: out_word = 8'hF5;
		16'hE2C1: out_word = 8'hCC;
		16'hE2C2: out_word = 8'hDC;
		16'hE2C3: out_word = 8'hD7;
		16'hE2C4: out_word = 8'h87;
		16'hE2C5: out_word = 8'hEF;
		16'hE2C6: out_word = 8'hDC;
		16'hE2C7: out_word = 8'h45;
		16'hE2C8: out_word = 8'h8F;
		16'hE2C9: out_word = 8'hEF;
		16'hE2CA: out_word = 8'hB9;
		16'hE2CB: out_word = 8'h07;
		16'hE2CC: out_word = 8'hEF;
		16'hE2CD: out_word = 8'hC3;
		16'hE2CE: out_word = 8'hFE;
		16'hE2CF: out_word = 8'h87;
		16'hE2D0: out_word = 8'hCD;
		16'hE2D1: out_word = 8'h18;
		16'hE2D2: out_word = 8'h8A;
		16'hE2D3: out_word = 8'hA7;
		16'hE2D4: out_word = 8'h20;
		16'hE2D5: out_word = 8'h08;
		16'hE2D6: out_word = 8'h17;
		16'hE2D7: out_word = 8'h6B;
		16'hE2D8: out_word = 8'h89;
		16'hE2D9: out_word = 8'h00;
		16'hE2DA: out_word = 8'h07;
		16'hE2DB: out_word = 8'hCC;
		16'hE2DC: out_word = 8'h9F;
		16'hE2DD: out_word = 8'h3A;
		16'hE2DE: out_word = 8'hF2;
		16'hE2DF: out_word = 8'h8A;
		16'hE2E0: out_word = 8'h8C;
		16'hE2E1: out_word = 8'h4C;
		16'hE2E2: out_word = 8'hF8;
		16'hE2E3: out_word = 8'hB1;
		16'hE2E4: out_word = 8'hF8;
		16'hE2E5: out_word = 8'h93;
		16'hE2E6: out_word = 8'h5E;
		16'hE2E7: out_word = 8'h37;
		16'hE2E8: out_word = 8'hC8;
		16'hE2E9: out_word = 8'h3D;
		16'hE2EA: out_word = 8'h11;
		16'hE2EB: out_word = 8'hB5;
		16'hE2EC: out_word = 8'hF8;
		16'hE2ED: out_word = 8'hD8;
		16'hE2EE: out_word = 8'h2A;
		16'hE2EF: out_word = 8'hF4;
		16'hE2F0: out_word = 8'hCF;
		16'hE2F1: out_word = 8'h23;
		16'hE2F2: out_word = 8'hFC;
		16'hE2F3: out_word = 8'h7E;
		16'hE2F4: out_word = 8'hED;
		16'hE2F5: out_word = 8'h5B;
		16'hE2F6: out_word = 8'hA7;
		16'hE2F7: out_word = 8'hB0;
		16'hE2F8: out_word = 8'hB1;
		16'hE2F9: out_word = 8'hA7;
		16'hE2FA: out_word = 8'hC9;
		16'hE2FB: out_word = 8'hDD;
		16'hE2FC: out_word = 8'hBB;
		16'hE2FD: out_word = 8'h7D;
		16'hE2FE: out_word = 8'h72;
		16'hE2FF: out_word = 8'hD8;
		16'hE300: out_word = 8'h1F;
		16'hE301: out_word = 8'hA1;
		16'hE302: out_word = 8'h89;
		16'hE303: out_word = 8'hF4;
		16'hE304: out_word = 8'hBF;
		16'hE305: out_word = 8'h3E;
		16'hE306: out_word = 8'hD7;
		16'hE307: out_word = 8'h05;
		16'hE308: out_word = 8'hF5;
		16'hE309: out_word = 8'h7A;
		16'hE30A: out_word = 8'h29;
		16'hE30B: out_word = 8'h42;
		16'hE30C: out_word = 8'h4B;
		16'hE30D: out_word = 8'hE5;
		16'hE30E: out_word = 8'h77;
		16'hE30F: out_word = 8'hBF;
		16'hE310: out_word = 8'h02;
		16'hE311: out_word = 8'h18;
		16'hE312: out_word = 8'h38;
		16'hE313: out_word = 8'h2D;
		16'hE314: out_word = 8'hEE;
		16'hE315: out_word = 8'h04;
		16'hE316: out_word = 8'h84;
		16'hE317: out_word = 8'hEE;
		16'hE318: out_word = 8'hB5;
		16'hE319: out_word = 8'hE0;
		16'hE31A: out_word = 8'hEE;
		16'hE31B: out_word = 8'h26;
		16'hE31C: out_word = 8'hF5;
		16'hE31D: out_word = 8'h7E;
		16'hE31E: out_word = 8'hCB;
		16'hE31F: out_word = 8'h7F;
		16'hE320: out_word = 8'h06;
		16'hE321: out_word = 8'hE0;
		16'hE322: out_word = 8'h28;
		16'hE323: out_word = 8'h02;
		16'hE324: out_word = 8'h25;
		16'hE325: out_word = 8'hF0;
		16'hE326: out_word = 8'h28;
		16'hE327: out_word = 8'hEA;
		16'hE328: out_word = 8'h4B;
		16'hE329: out_word = 8'h85;
		16'hE32A: out_word = 8'h6C;
		16'hE32B: out_word = 8'hEC;
		16'hE32C: out_word = 8'h12;
		16'hE32D: out_word = 8'hD1;
		16'hE32E: out_word = 8'hEC;
		16'hE32F: out_word = 8'h60;
		16'hE330: out_word = 8'h81;
		16'hE331: out_word = 8'h02;
		16'hE332: out_word = 8'hBE;
		16'hE333: out_word = 8'h91;
		16'hE334: out_word = 8'h01;
		16'hE335: out_word = 8'h43;
		16'hE336: out_word = 8'h8C;
		16'hE337: out_word = 8'h27;
		16'hE338: out_word = 8'h19;
		16'hE339: out_word = 8'h1C;
		16'hE33A: out_word = 8'h00;
		16'hE33B: out_word = 8'h04;
		16'hE33C: out_word = 8'h19;
		16'hE33D: out_word = 8'h7E;
		16'hE33E: out_word = 8'h7E;
		16'hE33F: out_word = 8'h85;
		16'hE340: out_word = 8'h28;
		16'hE341: out_word = 8'hFE;
		16'hE342: out_word = 8'hF5;
		16'hE343: out_word = 8'h80;
		16'hE344: out_word = 8'h20;
		16'hE345: out_word = 8'h09;
		16'hE346: out_word = 8'hFD;
		16'hE347: out_word = 8'h2C;
		16'hE348: out_word = 8'hDD;
		16'hE349: out_word = 8'h56;
		16'hE34A: out_word = 8'h89;
		16'hE34B: out_word = 8'h0D;
		16'hE34C: out_word = 8'h01;
		16'hE34D: out_word = 8'h0C;
		16'hE34E: out_word = 8'h72;
		16'hE34F: out_word = 8'hDB;
		16'hE350: out_word = 8'hFD;
		16'hE351: out_word = 8'hAB;
		16'hE352: out_word = 8'h00;
		16'hE353: out_word = 8'h79;
		16'hE354: out_word = 8'hFD;
		16'hE355: out_word = 8'hA7;
		16'hE356: out_word = 8'hE1;
		16'hE357: out_word = 8'hC2;
		16'hE358: out_word = 8'h8F;
		16'hE359: out_word = 8'h88;
		16'hE35A: out_word = 8'hE5;
		16'hE35B: out_word = 8'h3F;
		16'hE35C: out_word = 8'hD6;
		16'hE35D: out_word = 8'h4E;
		16'hE35E: out_word = 8'h0D;
		16'hE35F: out_word = 8'hAF;
		16'hE360: out_word = 8'h5F;
		16'hE361: out_word = 8'h06;
		16'hE362: out_word = 8'h08;
		16'hE363: out_word = 8'hCF;
		16'hE364: out_word = 8'hCB;
		16'hE365: out_word = 8'h19;
		16'hE366: out_word = 8'h04;
		16'hE367: out_word = 8'h10;
		16'hE368: out_word = 8'hFA;
		16'hE369: out_word = 8'h3D;
		16'hE36A: out_word = 8'h33;
		16'hE36B: out_word = 8'hDF;
		16'hE36C: out_word = 8'h1C;
		16'hE36D: out_word = 8'hD6;
		16'hE36E: out_word = 8'h0E;
		16'hE36F: out_word = 8'h17;
		16'hE370: out_word = 8'hB6;
		16'hE371: out_word = 8'h0F;
		16'hE372: out_word = 8'hB9;
		16'hE373: out_word = 8'h28;
		16'hE374: out_word = 8'hF7;
		16'hE375: out_word = 8'h13;
		16'hE376: out_word = 8'h37;
		16'hE377: out_word = 8'hF7;
		16'hE378: out_word = 8'h14;
		16'hE379: out_word = 8'h83;
		16'hE37A: out_word = 8'hEE;
		16'hE37B: out_word = 8'h33;
		16'hE37C: out_word = 8'hF7;
		16'hE37D: out_word = 8'h21;
		16'hE37E: out_word = 8'hFD;
		16'hE37F: out_word = 8'h22;
		16'hE380: out_word = 8'h47;
		16'hE381: out_word = 8'hFD;
		16'hE382: out_word = 8'hBC;
		16'hE383: out_word = 8'hF1;
		16'hE384: out_word = 8'h15;
		16'hE385: out_word = 8'hE6;
		16'hE386: out_word = 8'hF0;
		16'hE387: out_word = 8'hFE;
		16'hE388: out_word = 8'h64;
		16'hE389: out_word = 8'hF6;
		16'hE38A: out_word = 8'h85;
		16'hE38B: out_word = 8'h7B;
		16'hE38C: out_word = 8'h04;
		16'hE38D: out_word = 8'h8F;
		16'hE38E: out_word = 8'h33;
		16'hE38F: out_word = 8'hC0;
		16'hE390: out_word = 8'h8F;
		16'hE391: out_word = 8'h3B;
		16'hE392: out_word = 8'hF1;
		16'hE393: out_word = 8'h49;
		16'hE394: out_word = 8'h7C;
		16'hE395: out_word = 8'h00;
		16'hE396: out_word = 8'hCE;
		16'hE397: out_word = 8'hC1;
		16'hE398: out_word = 8'h04;
		16'hE399: out_word = 8'hE6;
		16'hE39A: out_word = 8'hAE;
		16'hE39B: out_word = 8'h4F;
		16'hE39C: out_word = 8'h78;
		16'hE39D: out_word = 8'h98;
		16'hE39E: out_word = 8'hAF;
		16'hE39F: out_word = 8'h71;
		16'hE3A0: out_word = 8'h23;
		16'hE3A1: out_word = 8'h70;
		16'hE3A2: out_word = 8'hD8;
		16'hE3A3: out_word = 8'h36;
		16'hE3A4: out_word = 8'hFF;
		16'hE3A5: out_word = 8'h76;
		16'hE3A6: out_word = 8'h77;
		16'hE3A7: out_word = 8'hCD;
		16'hE3A8: out_word = 8'hFE;
		16'hE3A9: out_word = 8'h11;
		16'hE3AA: out_word = 8'h08;
		16'hE3AB: out_word = 8'h51;
		16'hE3AC: out_word = 8'h60;
		16'hE3AD: out_word = 8'h7D;
		16'hE3AE: out_word = 8'hFA;
		16'hE3AF: out_word = 8'hDF;
		16'hE3B0: out_word = 8'hFC;
		16'hE3B1: out_word = 8'h5D;
		16'hE3B2: out_word = 8'h56;
		16'hE3B3: out_word = 8'h3E;
		16'hE3B4: out_word = 8'hF3;
		16'hE3B5: out_word = 8'h77;
		16'hE3B6: out_word = 8'hFA;
		16'hE3B7: out_word = 8'hC9;
		16'hE3B8: out_word = 8'hF1;
		16'hE3B9: out_word = 8'h9B;
		16'hE3BA: out_word = 8'h59;
		16'hE3BB: out_word = 8'h19;
		16'hE3BC: out_word = 8'hD9;
		16'hE3BD: out_word = 8'h21;
		16'hE3BE: out_word = 8'hC8;
		16'hE3BF: out_word = 8'hD9;
		16'hE3C0: out_word = 8'h26;
		16'hE3C1: out_word = 8'hF7;
		16'hE3C2: out_word = 8'h12;
		16'hE3C3: out_word = 8'h08;
		16'hE3C4: out_word = 8'h44;
		16'hE3C5: out_word = 8'h85;
		16'hE3C6: out_word = 8'h8B;
		16'hE3C7: out_word = 8'h09;
		16'hE3C8: out_word = 8'h0C;
		16'hE3C9: out_word = 8'h68;
		16'hE3CA: out_word = 8'h4D;
		16'hE3CB: out_word = 8'hCD;
		16'hE3CC: out_word = 8'h2F;
		16'hE3CD: out_word = 8'h7E;
		16'hE3CE: out_word = 8'hF8;
		16'hE3CF: out_word = 8'h2B;
		16'hE3D0: out_word = 8'hC5;
		16'hE3D1: out_word = 8'h4C;
		16'hE3D2: out_word = 8'hC9;
		16'hE3D3: out_word = 8'h43;
		16'hE3D4: out_word = 8'h71;
		16'hE3D5: out_word = 8'hCC;
		16'hE3D6: out_word = 8'hCE;
		16'hE3D7: out_word = 8'h70;
		16'hE3D8: out_word = 8'h01;
		16'hE3D9: out_word = 8'hF9;
		16'hE3DA: out_word = 8'h73;
		16'hE3DB: out_word = 8'h02;
		16'hE3DC: out_word = 8'h57;
		16'hE3DD: out_word = 8'hE0;
		16'hE3DE: out_word = 8'h26;
		16'hE3DF: out_word = 8'h25;
		16'hE3E0: out_word = 8'h13;
		16'hE3E1: out_word = 8'hFF;
		16'hE3E2: out_word = 8'h09;
		16'hE3E3: out_word = 8'hDB;
		16'hE3E4: out_word = 8'h9F;
		16'hE3E5: out_word = 8'h4B;
		16'hE3E6: out_word = 8'hDD;
		16'hE3E7: out_word = 8'h36;
		16'hE3E8: out_word = 8'h07;
		16'hE3E9: out_word = 8'h00;
		16'hE3EA: out_word = 8'h0E;
		16'hE3EB: out_word = 8'h85;
		16'hE3EC: out_word = 8'h08;
		16'hE3ED: out_word = 8'h09;
		16'hE3EE: out_word = 8'h40;
		16'hE3EF: out_word = 8'hC7;
		16'hE3F0: out_word = 8'h8D;
		16'hE3F1: out_word = 8'h42;
		16'hE3F2: out_word = 8'hBE;
		16'hE3F3: out_word = 8'hA7;
		16'hE3F4: out_word = 8'hFF;
		16'hE3F5: out_word = 8'h94;
		16'hE3F6: out_word = 8'h21;
		16'hE3F7: out_word = 8'hF2;
		16'hE3F8: out_word = 8'hCF;
		16'hE3F9: out_word = 8'hBE;
		16'hE3FA: out_word = 8'h3F;
		16'hE3FB: out_word = 8'hD8;
		16'hE3FC: out_word = 8'hC2;
		16'hE3FD: out_word = 8'h32;
		16'hE3FE: out_word = 8'hF3;
		16'hE3FF: out_word = 8'h69;
		16'hE400: out_word = 8'h88;
		16'hE401: out_word = 8'h2A;
		16'hE402: out_word = 8'h11;
		16'hE403: out_word = 8'h7E;
		16'hE404: out_word = 8'hCF;
		16'hE405: out_word = 8'h19;
		16'hE406: out_word = 8'h22;
		16'hE407: out_word = 8'hF4;
		16'hE408: out_word = 8'h24;
		16'hE409: out_word = 8'h7E;
		16'hE40A: out_word = 8'hF1;
		16'hE40B: out_word = 8'h52;
		16'hE40C: out_word = 8'h38;
		16'hE40D: out_word = 8'h16;
		16'hE40E: out_word = 8'hD6;
		16'hE40F: out_word = 8'h3E;
		16'hE410: out_word = 8'h21;
		16'hE411: out_word = 8'h8A;
		16'hE412: out_word = 8'h8C;
		16'hE413: out_word = 8'h28;
		16'hE414: out_word = 8'h0F;
		16'hE415: out_word = 8'h70;
		16'hE416: out_word = 8'hDD;
		16'hE417: out_word = 8'h6B;
		16'hE418: out_word = 8'h89;
		16'hE419: out_word = 8'hA6;
		16'hE41A: out_word = 8'h09;
		16'hE41B: out_word = 8'hFA;
		16'hE41C: out_word = 8'h22;
		16'hE41D: out_word = 8'h61;
		16'hE41E: out_word = 8'hFA;
		16'hE41F: out_word = 8'h03;
		16'hE420: out_word = 8'hC3;
		16'hE421: out_word = 8'h3C;
		16'hE422: out_word = 8'h07;
		16'hE423: out_word = 8'hF0;
		16'hE424: out_word = 8'hCF;
		16'hE425: out_word = 8'hFF;
		16'hE426: out_word = 8'hAF;
		16'hE427: out_word = 8'hC9;
		16'hE428: out_word = 8'hF5;
		16'hE429: out_word = 8'hE5;
		16'hE42A: out_word = 8'h78;
		16'hE42B: out_word = 8'hE6;
		16'hE42C: out_word = 8'h0F;
		16'hE42D: out_word = 8'h47;
		16'hE42E: out_word = 8'h77;
		16'hE42F: out_word = 8'hE0;
		16'hE430: out_word = 8'h5C;
		16'hE431: out_word = 8'h7E;
		16'hE432: out_word = 8'h5D;
		16'hE433: out_word = 8'h01;
		16'hE434: out_word = 8'h4F;
		16'hE435: out_word = 8'hE1;
		16'hE436: out_word = 8'hF6;
		16'hE437: out_word = 8'hE0;
		16'hE438: out_word = 8'hB0;
		16'hE439: out_word = 8'h47;
		16'hE43A: out_word = 8'hFB;
		16'hE43B: out_word = 8'hE1;
		16'hE43C: out_word = 8'hF1;
		16'hE43D: out_word = 8'hC3;
		16'hE43E: out_word = 8'h12;
		16'hE43F: out_word = 8'h8E;
		16'hE440: out_word = 8'h16;
		16'hE441: out_word = 8'h7F;
		16'hE442: out_word = 8'hE6;
		16'hE443: out_word = 8'h45;
		16'hE444: out_word = 8'h8F;
		16'hE445: out_word = 8'hFE;
		16'hE446: out_word = 8'h06;
		16'hE447: out_word = 8'h1E;
		16'hE448: out_word = 8'h01;
		16'hE449: out_word = 8'hC8;
		16'hE44A: out_word = 8'h0E;
		16'hE44B: out_word = 8'h0E;
		16'hE44C: out_word = 8'h60;
		16'hE44D: out_word = 8'hFD;
		16'hE44E: out_word = 8'h0B;
		16'hE44F: out_word = 8'h4C;
		16'hE450: out_word = 8'h02;
		16'hE451: out_word = 8'hFB;
		16'hE452: out_word = 8'h0C;
		16'hE453: out_word = 8'hC0;
		16'hE454: out_word = 8'hFD;
		16'hE455: out_word = 8'h01;
		16'hE456: out_word = 8'hB5;
		16'hE457: out_word = 8'h00;
		16'hE458: out_word = 8'hF7;
		16'hE459: out_word = 8'hA4;
		16'hE45A: out_word = 8'hE5;
		16'hE45B: out_word = 8'h21;
		16'hE45C: out_word = 8'h82;
		16'hE45D: out_word = 8'hFD;
		16'hE45E: out_word = 8'h89;
		16'hE45F: out_word = 8'h85;
		16'hE460: out_word = 8'h6F;
		16'hE461: out_word = 8'h3E;
		16'hE462: out_word = 8'h00;
		16'hE463: out_word = 8'h8C;
		16'hE464: out_word = 8'hB7;
		16'hE465: out_word = 8'hB8;
		16'hE466: out_word = 8'hAD;
		16'hE467: out_word = 8'hC5;
		16'hE468: out_word = 8'h89;
		16'hE469: out_word = 8'hC1;
		16'hE46A: out_word = 8'hD1;
		16'hE46B: out_word = 8'h8F;
		16'hE46C: out_word = 8'h21;
		16'hE46D: out_word = 8'h8A;
		16'hE46E: out_word = 8'h7C;
		16'hE46F: out_word = 8'h08;
		16'hE470: out_word = 8'h3E;
		16'hE471: out_word = 8'h03;
		16'hE472: out_word = 8'h18;
		16'hE473: out_word = 8'h05;
		16'hE474: out_word = 8'h49;
		16'hE475: out_word = 8'h01;
		16'hE476: out_word = 8'hF9;
		16'hE477: out_word = 8'hE7;
		16'hE478: out_word = 8'h02;
		16'hE479: out_word = 8'hCD;
		16'hE47A: out_word = 8'hD7;
		16'hE47B: out_word = 8'hF3;
		16'hE47C: out_word = 8'hD5;
		16'hE47D: out_word = 8'hC5;
		16'hE47E: out_word = 8'hE1;
		16'hE47F: out_word = 8'h01;
		16'hE480: out_word = 8'hB3;
		16'hE481: out_word = 8'h00;
		16'hE482: out_word = 8'h7C;
		16'hE483: out_word = 8'hD3;
		16'hE484: out_word = 8'hBB;
		16'hE485: out_word = 8'hCD;
		16'hE486: out_word = 8'h12;
		16'hE487: out_word = 8'h8A;
		16'hE488: out_word = 8'h98;
		16'hE489: out_word = 8'h58;
		16'hE48A: out_word = 8'hEE;
		16'hE48B: out_word = 8'h0C;
		16'hE48C: out_word = 8'h5F;
		16'hE48D: out_word = 8'hED;
		16'hE48E: out_word = 8'hA2;
		16'hE48F: out_word = 8'h1B;
		16'hE490: out_word = 8'h7A;
		16'hE491: out_word = 8'hB3;
		16'hE492: out_word = 8'hD2;
		16'hE493: out_word = 8'h20;
		16'hE494: out_word = 8'hF6;
		16'hE495: out_word = 8'h32;
		16'hE496: out_word = 8'hE9;
		16'hE497: out_word = 8'hE7;
		16'hE498: out_word = 8'hF2;
		16'hE499: out_word = 8'h78;
		16'hE49A: out_word = 8'hFE;
		16'hE49B: out_word = 8'h77;
		16'hE49C: out_word = 8'hF2;
		16'hE49D: out_word = 8'h20;
		16'hE49E: out_word = 8'hFA;
		16'hE49F: out_word = 8'hC1;
		16'hE4A0: out_word = 8'hD1;
		16'hE4A1: out_word = 8'h61;
		16'hE4A2: out_word = 8'h63;
		16'hE4A3: out_word = 8'hCE;
		16'hE4A4: out_word = 8'h18;
		16'hE4A5: out_word = 8'h04;
		16'hE4A6: out_word = 8'h89;
		16'hE4A7: out_word = 8'hCE;
		16'hE4A8: out_word = 8'hEB;
		16'hE4A9: out_word = 8'hDB;
		16'hE4AA: out_word = 8'hA5;
		16'hE4AB: out_word = 8'hB3;
		16'hE4AC: out_word = 8'hEB;
		16'hE4AD: out_word = 8'h02;
		16'hE4AE: out_word = 8'hC1;
		16'hE4AF: out_word = 8'hED;
		16'hE4B0: out_word = 8'h70;
		16'hE4B1: out_word = 8'hD3;
		16'hE4B2: out_word = 8'hB3;
		16'hE4B3: out_word = 8'hEF;
		16'hE4B4: out_word = 8'h1E;
		16'hE4B5: out_word = 8'h48;
		16'hE4B6: out_word = 8'hC3;
		16'hE4B7: out_word = 8'h78;
		16'hE4B8: out_word = 8'hF6;
		16'hE4B9: out_word = 8'h50;
		16'hE4BA: out_word = 8'h06;
		16'hE4BB: out_word = 8'hAF;
		16'hE4BC: out_word = 8'h79;
		16'hE4BD: out_word = 8'h5E;
		16'hE4BE: out_word = 8'hFA;
		16'hE4BF: out_word = 8'h7A;
		16'hE4C0: out_word = 8'hFA;
		16'hE4C1: out_word = 8'hBC;
		16'hE4C2: out_word = 8'h7B;
		16'hE4C3: out_word = 8'hFA;
		16'hE4C4: out_word = 8'h42;
		16'hE4C5: out_word = 8'hA5;
		16'hE4C6: out_word = 8'h15;
		16'hE4C7: out_word = 8'hBC;
		16'hE4C8: out_word = 8'h3F;
		16'hE4C9: out_word = 8'h7F;
		16'hE4CA: out_word = 8'hC9;
		16'hE4CB: out_word = 8'hDB;
		16'hE4CC: out_word = 8'hBB;
		16'hE4CD: out_word = 8'h17;
		16'hE4CE: out_word = 8'h38;
		16'hE4CF: out_word = 8'hFB;
		16'hE4D0: out_word = 8'h72;
		16'hE4D1: out_word = 8'hFA;
		16'hE4D2: out_word = 8'h30;
		16'hE4D3: out_word = 8'hE5;
		16'hE4D4: out_word = 8'hFA;
		16'hE4D5: out_word = 8'h1F;
		16'hE4D6: out_word = 8'h3C;
		16'hE4D7: out_word = 8'hF4;
		16'hE4D8: out_word = 8'h3E;
		16'hE4D9: out_word = 8'h80;
		16'hE4DA: out_word = 8'hD3;
		16'hE4DB: out_word = 8'h33;
		16'hE4DC: out_word = 8'h28;
		16'hE4DD: out_word = 8'h76;
		16'hE4DE: out_word = 8'hF0;
		16'hE4DF: out_word = 8'hF3;
		16'hE4E0: out_word = 8'h06;
		16'hE4E1: out_word = 8'hC9;
		16'hE4E2: out_word = 8'h06;
		16'hE4E3: out_word = 8'h30;
		16'hE4E4: out_word = 8'hB7;
		16'hE4E5: out_word = 8'hF6;
		16'hE4E6: out_word = 8'h07;
		16'hE4E7: out_word = 8'h05;
		16'hE4E8: out_word = 8'h28;
		16'hE4E9: out_word = 8'hB9;
		16'hE4EA: out_word = 8'hA8;
		16'hE4EB: out_word = 8'hE6;
		16'hE4EC: out_word = 8'hF5;
		16'hE4ED: out_word = 8'h42;
		16'hE4EE: out_word = 8'h69;
		16'hE4EF: out_word = 8'h83;
		16'hE4F0: out_word = 8'h70;
		16'hE4F1: out_word = 8'h6D;
		16'hE4F2: out_word = 8'h03;
		16'hE4F3: out_word = 8'h21;
		16'hE4F4: out_word = 8'h60;
		16'hE4F5: out_word = 8'h5B;
		16'hE4F6: out_word = 8'h77;
		16'hE4F7: out_word = 8'h59;
		16'hE4F8: out_word = 8'h3E;
		16'hE4F9: out_word = 8'h14;
		16'hE4FA: out_word = 8'hB4;
		16'hE4FB: out_word = 8'h9B;
		16'hE4FC: out_word = 8'hED;
		16'hE4FD: out_word = 8'h51;
		16'hE4FE: out_word = 8'hAE;
		16'hE4FF: out_word = 8'h0E;
		16'hE500: out_word = 8'h69;
		16'hE501: out_word = 8'hE5;
		16'hE502: out_word = 8'hFB;
		16'hE503: out_word = 8'h61;
		16'hE504: out_word = 8'h09;
		16'hE505: out_word = 8'hFB;
		16'hE506: out_word = 8'h1E;
		16'hE507: out_word = 8'hF8;
		16'hE508: out_word = 8'hA3;
		16'hE509: out_word = 8'hA3;
		16'hE50A: out_word = 8'hF8;
		16'hE50B: out_word = 8'hC8;
		16'hE50C: out_word = 8'h4F;
		16'hE50D: out_word = 8'hD8;
		16'hE50E: out_word = 8'hB1;
		16'hE50F: out_word = 8'hBE;
		16'hE510: out_word = 8'h13;
		16'hE511: out_word = 8'h78;
		16'hE512: out_word = 8'hD8;
		16'hE513: out_word = 8'hA1;
		16'hE514: out_word = 8'hE2;
		16'hE515: out_word = 8'hAD;
		16'hE516: out_word = 8'hAF;
		16'hE517: out_word = 8'h9F;
		16'hE518: out_word = 8'h03;
		16'hE519: out_word = 8'h57;
		16'hE51A: out_word = 8'h05;
		16'hE51B: out_word = 8'hCA;
		16'hE51C: out_word = 8'hD4;
		16'hE51D: out_word = 8'h89;
		16'hE51E: out_word = 8'h32;
		16'hE51F: out_word = 8'h53;
		16'hE520: out_word = 8'hC2;
		16'hE521: out_word = 8'hFB;
		16'hE522: out_word = 8'h4F;
		16'hE523: out_word = 8'h52;
		16'hE524: out_word = 8'h9D;
		16'hE525: out_word = 8'h9C;
		16'hE526: out_word = 8'hD3;
		16'hE527: out_word = 8'h11;
		16'hE528: out_word = 8'hF0;
		16'hE529: out_word = 8'hCD;
		16'hE52A: out_word = 8'h35;
		16'hE52B: out_word = 8'h5B;
		16'hE52C: out_word = 8'hA7;
		16'hE52D: out_word = 8'h2A;
		16'hE52E: out_word = 8'h77;
		16'hE52F: out_word = 8'h9C;
		16'hE530: out_word = 8'h29;
		16'hE531: out_word = 8'hCC;
		16'hE532: out_word = 8'hD3;
		16'hE533: out_word = 8'h03;
		16'hE534: out_word = 8'h6F;
		16'hE535: out_word = 8'h05;
		16'hE536: out_word = 8'hC2;
		16'hE537: out_word = 8'h6E;
		16'hE538: out_word = 8'h02;
		16'hE539: out_word = 8'hFC;
		16'hE53A: out_word = 8'hF3;
		16'hE53B: out_word = 8'hDB;
		16'hE53C: out_word = 8'h0F;
		16'hE53D: out_word = 8'hCB;
		16'hE53E: out_word = 8'h8F;
		16'hE53F: out_word = 8'hD3;
		16'hE540: out_word = 8'h43;
		16'hE541: out_word = 8'hC2;
		16'hE542: out_word = 8'h1D;
		16'hE543: out_word = 8'hFF;
		16'hE544: out_word = 8'h22;
		16'hE545: out_word = 8'h3C;
		16'hE546: out_word = 8'h03;
		16'hE547: out_word = 8'h11;
		16'hE548: out_word = 8'h44;
		16'hE549: out_word = 8'h5B;
		16'hE54A: out_word = 8'h01;
		16'hE54B: out_word = 8'hC4;
		16'hE54C: out_word = 8'h1B;
		16'hE54D: out_word = 8'hEB;
		16'hE54E: out_word = 8'hED;
		16'hE54F: out_word = 8'hA4;
		16'hE550: out_word = 8'hB0;
		16'hE551: out_word = 8'hEB;
		16'hE552: out_word = 8'hCF;
		16'hE553: out_word = 8'hC9;
		16'hE554: out_word = 8'hEB;
		16'hE555: out_word = 8'hC3;
		16'hE556: out_word = 8'hE1;
		16'hE557: out_word = 8'hF7;
		16'hE558: out_word = 8'hA4;
		16'hE559: out_word = 8'hE6;
		16'hE55A: out_word = 8'hF7;
		16'hE55B: out_word = 8'h57;
		16'hE55C: out_word = 8'hFE;
		16'hE55D: out_word = 8'hF9;
		16'hE55E: out_word = 8'hBA;
		16'hE55F: out_word = 8'h3E;
		16'hE560: out_word = 8'h00;
		16'hE561: out_word = 8'hC8;
		16'hE562: out_word = 8'h3D;
		16'hE563: out_word = 8'hC9;
		16'hE564: out_word = 8'h66;
		16'hE565: out_word = 8'hD2;
		16'hE566: out_word = 8'h02;
		16'hE567: out_word = 8'hCA;
		16'hE568: out_word = 8'h21;
		16'hE569: out_word = 8'h7E;
		16'hE56A: out_word = 8'hE9;
		16'hE56B: out_word = 8'hE5;
		16'hE56C: out_word = 8'h87;
		16'hE56D: out_word = 8'h5F;
		16'hE56E: out_word = 8'h16;
		16'hE56F: out_word = 8'h00;
		16'hE570: out_word = 8'h06;
		16'hE571: out_word = 8'h33;
		16'hE572: out_word = 8'h1D;
		16'hE573: out_word = 8'hF8;
		16'hE574: out_word = 8'h73;
		16'hE575: out_word = 8'hC2;
		16'hE576: out_word = 8'hCD;
		16'hE577: out_word = 8'hBE;
		16'hE578: out_word = 8'h1E;
		16'hE579: out_word = 8'hE9;
		16'hE57A: out_word = 8'h47;
		16'hE57B: out_word = 8'h7A;
		16'hE57C: out_word = 8'hFA;
		16'hE57D: out_word = 8'h4F;
		16'hE57E: out_word = 8'hF5;
		16'hE57F: out_word = 8'hFA;
		16'hE580: out_word = 8'h57;
		16'hE581: out_word = 8'hEB;
		16'hE582: out_word = 8'hFA;
		16'hE583: out_word = 8'h5F;
		16'hE584: out_word = 8'hDE;
		16'hE585: out_word = 8'hFA;
		16'hE586: out_word = 8'hE9;
		16'hE587: out_word = 8'h43;
		16'hE588: out_word = 8'h1D;
		16'hE589: out_word = 8'hC0;
		16'hE58A: out_word = 8'h37;
		16'hE58B: out_word = 8'h79;
		16'hE58C: out_word = 8'h1E;
		16'hE58D: out_word = 8'h90;
		16'hE58E: out_word = 8'h1B;
		16'hE58F: out_word = 8'hCD;
		16'hE590: out_word = 8'hC3;
		16'hE591: out_word = 8'h07;
		16'hE592: out_word = 8'h3E;
		16'hE593: out_word = 8'hEE;
		16'hE594: out_word = 8'h12;
		16'hE595: out_word = 8'hB6;
		16'hE596: out_word = 8'hE7;
		16'hE597: out_word = 8'hF8;
		16'hE598: out_word = 8'h01;
		16'hE599: out_word = 8'h13;
		16'hE59A: out_word = 8'h00;
		16'hE59B: out_word = 8'hE6;
		16'hE59C: out_word = 8'h11;
		16'hE59D: out_word = 8'hFF;
		16'hE59E: out_word = 8'h20;
		16'hE59F: out_word = 8'h2A;
		16'hE5A0: out_word = 8'h15;
		16'hE5A1: out_word = 8'h27;
		16'hE5A2: out_word = 8'hFB;
		16'hE5A3: out_word = 8'h01;
		16'hE5A4: out_word = 8'h14;
		16'hE5A5: out_word = 8'hF9;
		16'hE5A6: out_word = 8'h00;
		16'hE5A7: out_word = 8'hAF;
		16'hE5A8: out_word = 8'h08;
		16'hE5A9: out_word = 8'h21;
		16'hE5AA: out_word = 8'h48;
		16'hE5AB: out_word = 8'hEA;
		16'hE5AC: out_word = 8'hC5;
		16'hE5AD: out_word = 8'hD1;
		16'hE5AE: out_word = 8'h1D;
		16'hE5AF: out_word = 8'h85;
		16'hE5B0: out_word = 8'h3A;
		16'hE5B1: out_word = 8'h08;
		16'hE5B2: out_word = 8'hEB;
		16'hE5B3: out_word = 8'h3D;
		16'hE5B4: out_word = 8'h28;
		16'hE5B5: out_word = 8'hD8;
		16'hE5B6: out_word = 8'hFD;
		16'hE5B7: out_word = 8'h87;
		16'hE5B8: out_word = 8'hEF;
		16'hE5B9: out_word = 8'h21;
		16'hE5BA: out_word = 8'h4E;
		16'hE5BB: out_word = 8'hAB;
		16'hE5BC: out_word = 8'hEF;
		16'hE5BD: out_word = 8'hED;
		16'hE5BE: out_word = 8'h60;
		16'hE5BF: out_word = 8'hB6;
		16'hE5C0: out_word = 8'h00;
		16'hE5C1: out_word = 8'h2E;
		16'hE5C2: out_word = 8'hFD;
		16'hE5C3: out_word = 8'h7E;
		16'hE5C4: out_word = 8'hAB;
		16'hE5C5: out_word = 8'hCB;
		16'hE5C6: out_word = 8'h57;
		16'hE5C7: out_word = 8'h20;
		16'hE5C8: out_word = 8'h02;
		16'hE5C9: out_word = 8'h26;
		16'hE5CA: out_word = 8'h40;
		16'hE5CB: out_word = 8'h77;
		16'hE5CC: out_word = 8'h41;
		16'hE5CD: out_word = 8'hCD;
		16'hE5CE: out_word = 8'hDC;
		16'hE5CF: out_word = 8'h13;
		16'hE5D0: out_word = 8'hE4;
		16'hE5D1: out_word = 8'hBA;
		16'hE5D2: out_word = 8'h3E;
		16'hE5D3: out_word = 8'h69;
		16'hE5D4: out_word = 8'hC3;
		16'hE5D5: out_word = 8'hED;
		16'hE5D6: out_word = 8'h79;
		16'hE5D7: out_word = 8'h20;
		16'hE5D8: out_word = 8'h13;
		16'hE5D9: out_word = 8'h17;
		16'hE5DA: out_word = 8'h07;
		16'hE5DB: out_word = 8'h8C;
		16'hE5DC: out_word = 8'hFD;
		16'hE5DD: out_word = 8'h01;
		16'hE5DE: out_word = 8'hFF;
		16'hE5DF: out_word = 8'hA7;
		16'hE5E0: out_word = 8'hF0;
		16'hE5E1: out_word = 8'hE6;
		16'hE5E2: out_word = 8'hA7;
		16'hE5E3: out_word = 8'h20;
		16'hE5E4: out_word = 8'hDB;
		16'hE5E5: out_word = 8'hD1;
		16'hE5E6: out_word = 8'h3E;
		16'hE5E7: out_word = 8'h7B;
		16'hE5E8: out_word = 8'hDB;
		16'hE5E9: out_word = 8'hEE;
		16'hE5EA: out_word = 8'hF5;
		16'hE5EB: out_word = 8'hF5;
		16'hE5EC: out_word = 8'h21;
		16'hE5ED: out_word = 8'h54;
		16'hE5EE: out_word = 8'hD4;
		16'hE5EF: out_word = 8'hB3;
		16'hE5F0: out_word = 8'h78;
		16'hE5F1: out_word = 8'hF4;
		16'hE5F2: out_word = 8'hF4;
		16'hE5F3: out_word = 8'hC3;
		16'hE5F4: out_word = 8'hB1;
		16'hE5F5: out_word = 8'h5F;
		16'hE5F6: out_word = 8'hF5;
		16'hE5F7: out_word = 8'h3E;
		16'hE5F8: out_word = 8'h81;
		16'hE5F9: out_word = 8'hD3;
		16'hE5FA: out_word = 8'h11;
		16'hE5FB: out_word = 8'h5C;
		16'hE5FC: out_word = 8'h1B;
		16'hE5FD: out_word = 8'h06;
		16'hE5FE: out_word = 8'h01;
		16'hE5FF: out_word = 8'hE7;
		16'hE600: out_word = 8'hF9;
		16'hE601: out_word = 8'hCD;
		16'hE602: out_word = 8'hCA;
		16'hE603: out_word = 8'h1D;
		16'hE604: out_word = 8'h9E;
		16'hE605: out_word = 8'hC5;
		16'hE606: out_word = 8'hB7;
		16'hE607: out_word = 8'h06;
		16'hE608: out_word = 8'hED;
		16'hE609: out_word = 8'hB3;
		16'hE60A: out_word = 8'hA2;
		16'hE60B: out_word = 8'h71;
		16'hE60C: out_word = 8'h88;
		16'hE60D: out_word = 8'hF4;
		16'hE60E: out_word = 8'hAC;
		16'hE60F: out_word = 8'h68;
		16'hE610: out_word = 8'hBE;
		16'hE611: out_word = 8'hAF;
		16'hE612: out_word = 8'hAB;
		16'hE613: out_word = 8'hD9;
		16'hE614: out_word = 8'hFD;
		16'hE615: out_word = 8'h3D;
		16'hE616: out_word = 8'h57;
		16'hE617: out_word = 8'h70;
		16'hE618: out_word = 8'h55;
		16'hE619: out_word = 8'h8F;
		16'hE61A: out_word = 8'hC6;
		16'hE61B: out_word = 8'hC5;
		16'hE61C: out_word = 8'hF5;
		16'hE61D: out_word = 8'hD0;
		16'hE61E: out_word = 8'h3E;
		16'hE61F: out_word = 8'h7A;
		16'hE620: out_word = 8'h54;
		16'hE621: out_word = 8'hBD;
		16'hE622: out_word = 8'hAB;
		16'hE623: out_word = 8'h6A;
		16'hE624: out_word = 8'h78;
		16'hE625: out_word = 8'h6E;
		16'hE626: out_word = 8'h6A;
		16'hE627: out_word = 8'hFE;
		16'hE628: out_word = 8'hCB;
		16'hE629: out_word = 8'h77;
		16'hE62A: out_word = 8'hE1;
		16'hE62B: out_word = 8'h20;
		16'hE62C: out_word = 8'h0A;
		16'hE62D: out_word = 8'hEB;
		16'hE62E: out_word = 8'h29;
		16'hE62F: out_word = 8'h37;
		16'hE630: out_word = 8'hED;
		16'hE631: out_word = 8'h6A;
		16'hE632: out_word = 8'h65;
		16'hE633: out_word = 8'h1B;
		16'hE634: out_word = 8'h53;
		16'hE635: out_word = 8'h1E;
		16'hE636: out_word = 8'hD1;
		16'hE637: out_word = 8'h00;
		16'hE638: out_word = 8'hF1;
		16'hE639: out_word = 8'hBF;
		16'hE63A: out_word = 8'h90;
		16'hE63B: out_word = 8'h6D;
		16'hE63C: out_word = 8'h84;
		16'hE63D: out_word = 8'h51;
		16'hE63E: out_word = 8'h4A;
		16'hE63F: out_word = 8'h1C;
		16'hE640: out_word = 8'h6D;
		16'hE641: out_word = 8'h29;
		16'hE642: out_word = 8'hBE;
		16'hE643: out_word = 8'hD3;
		16'hE644: out_word = 8'h7E;
		16'hE645: out_word = 8'hD5;
		16'hE646: out_word = 8'h0E;
		16'hE647: out_word = 8'hDB;
		16'hE648: out_word = 8'h14;
		16'hE649: out_word = 8'h89;
		16'hE64A: out_word = 8'hBB;
		16'hE64B: out_word = 8'h03;
		16'hE64C: out_word = 8'h3E;
		16'hE64D: out_word = 8'h0B;
		16'hE64E: out_word = 8'hF8;
		16'hE64F: out_word = 8'hD1;
		16'hE650: out_word = 8'hC9;
		16'hE651: out_word = 8'h40;
		16'hE652: out_word = 8'hEF;
		16'hE653: out_word = 8'h6B;
		16'hE654: out_word = 8'hF2;
		16'hE655: out_word = 8'h95;
		16'hE656: out_word = 8'h48;
		16'hE657: out_word = 8'h1C;
		16'hE658: out_word = 8'hBA;
		16'hE659: out_word = 8'hAA;
		16'hE65A: out_word = 8'h87;
		16'hE65B: out_word = 8'h50;
		16'hE65C: out_word = 8'hC0;
		16'hE65D: out_word = 8'hFA;
		16'hE65E: out_word = 8'h02;
		16'hE65F: out_word = 8'hFF;
		16'hE660: out_word = 8'hFF;
		16'hE661: out_word = 8'hDB;
		16'hE662: out_word = 8'h04;
		16'hE663: out_word = 8'h1F;
		16'hE664: out_word = 8'h30;
		16'hE665: out_word = 8'hFB;
		16'hE666: out_word = 8'hD3;
		16'hE667: out_word = 8'h05;
		16'hE668: out_word = 8'h49;
		16'hE669: out_word = 8'h9C;
		16'hE66A: out_word = 8'h21;
		16'hE66B: out_word = 8'hF1;
		16'hE66C: out_word = 8'h3F;
		16'hE66D: out_word = 8'h9F;
		16'hE66E: out_word = 8'h2B;
		16'hE66F: out_word = 8'hD3;
		16'hE670: out_word = 8'h03;
		16'hE671: out_word = 8'hCD;
		16'hE672: out_word = 8'hB8;
		16'hE673: out_word = 8'hE5;
		16'hE674: out_word = 8'h1E;
		16'hE675: out_word = 8'h7C;
		16'hE676: out_word = 8'hB5;
		16'hE677: out_word = 8'h4D;
		16'hE678: out_word = 8'hC1;
		16'hE679: out_word = 8'h93;
		16'hE67A: out_word = 8'h7E;
		16'hE67B: out_word = 8'hC9;
		16'hE67C: out_word = 8'h3E;
		16'hE67D: out_word = 8'h51;
		16'hE67E: out_word = 8'hCD;
		16'hE67F: out_word = 8'hF6;
		16'hE680: out_word = 8'hE4;
		16'hE681: out_word = 8'h85;
		16'hE682: out_word = 8'hFE;
		16'hE683: out_word = 8'h7C;
		16'hE684: out_word = 8'h20;
		16'hE685: out_word = 8'hF9;
		16'hE686: out_word = 8'h18;
		16'hE687: out_word = 8'h5A;
		16'hE688: out_word = 8'h29;
		16'hE689: out_word = 8'hF6;
		16'hE68A: out_word = 8'h3C;
		16'hE68B: out_word = 8'hFE;
		16'hE68C: out_word = 8'h20;
		16'hE68D: out_word = 8'hFA;
		16'hE68E: out_word = 8'h18;
		16'hE68F: out_word = 8'h21;
		16'hE690: out_word = 8'h08;
		16'hE691: out_word = 8'h3E;
		16'hE692: out_word = 8'h52;
		16'hE693: out_word = 8'h81;
		16'hE694: out_word = 8'hE8;
		16'hE695: out_word = 8'h02;
		16'hE696: out_word = 8'hC8;
		16'hE697: out_word = 8'h2F;
		16'hE698: out_word = 8'hE6;
		16'hE699: out_word = 8'hF4;
		16'hE69A: out_word = 8'hC1;
		16'hE69B: out_word = 8'hF1;
		16'hE69C: out_word = 8'h3E;
		16'hE69D: out_word = 8'h4C;
		16'hE69E: out_word = 8'h58;
		16'hE69F: out_word = 8'h68;
		16'hE6A0: out_word = 8'hDD;
		16'hE6A1: out_word = 8'h77;
		16'hE6A2: out_word = 8'hE4;
		16'hE6A3: out_word = 8'h8A;
		16'hE6A4: out_word = 8'h77;
		16'hE6A5: out_word = 8'hB4;
		16'hE6A6: out_word = 8'hBF;
		16'hE6A7: out_word = 8'hA2;
		16'hE6A8: out_word = 8'hC1;
		16'hE6A9: out_word = 8'h88;
		16'hE6AA: out_word = 8'h2F;
		16'hE6AB: out_word = 8'h37;
		16'hE6AC: out_word = 8'h88;
		16'hE6AD: out_word = 8'hEE;
		16'hE6AE: out_word = 8'hE1;
		16'hE6AF: out_word = 8'hA1;
		16'hE6B0: out_word = 8'h8C;
		16'hE6B1: out_word = 8'hCB;
		16'hE6B2: out_word = 8'hDF;
		16'hE6B3: out_word = 8'h8E;
		16'hE6B4: out_word = 8'hA9;
		16'hE6B5: out_word = 8'h8C;
		16'hE6B6: out_word = 8'h2F;
		16'hE6B7: out_word = 8'hC6;
		16'hE6B8: out_word = 8'h8D;
		16'hE6B9: out_word = 8'hFA;
		16'hE6BA: out_word = 8'h89;
		16'hE6BB: out_word = 8'hD6;
		16'hE6BC: out_word = 8'hCD;
		16'hE6BD: out_word = 8'h83;
		16'hE6BE: out_word = 8'h20;
		16'hE6BF: out_word = 8'h01;
		16'hE6C0: out_word = 8'hAF;
		16'hE6C1: out_word = 8'h57;
		16'hE6C2: out_word = 8'hDF;
		16'hE6C3: out_word = 8'h60;
		16'hE6C4: out_word = 8'h10;
		16'hE6C5: out_word = 8'hF5;
		16'hE6C6: out_word = 8'h60;
		16'hE6C7: out_word = 8'hF9;
		16'hE6C8: out_word = 8'h63;
		16'hE6C9: out_word = 8'hB3;
		16'hE6CA: out_word = 8'hED;
		16'hE6CB: out_word = 8'h98;
		16'hE6CC: out_word = 8'h3C;
		16'hE6CD: out_word = 8'hFD;
		16'hE6CE: out_word = 8'hA5;
		16'hE6CF: out_word = 8'h4B;
		16'hE6D0: out_word = 8'hF7;
		16'hE6D1: out_word = 8'h63;
		16'hE6D2: out_word = 8'h64;
		16'hE6D3: out_word = 8'hFE;
		16'hE6D4: out_word = 8'h63;
		16'hE6D5: out_word = 8'hB9;
		16'hE6D6: out_word = 8'hD4;
		16'hE6D7: out_word = 8'hEF;
		16'hE6D8: out_word = 8'hC5;
		16'hE6D9: out_word = 8'h7F;
		16'hE6DA: out_word = 8'h63;
		16'hE6DB: out_word = 8'h47;
		16'hE6DC: out_word = 8'h71;
		16'hE6DD: out_word = 8'hE4;
		16'hE6DE: out_word = 8'h89;
		16'hE6DF: out_word = 8'hFC;
		16'hE6E0: out_word = 8'h66;
		16'hE6E1: out_word = 8'hF5;
		16'hE6E2: out_word = 8'hE9;
		16'hE6E3: out_word = 8'hA7;
		16'hE6E4: out_word = 8'h20;
		16'hE6E5: out_word = 8'hDE;
		16'hE6E6: out_word = 8'hF7;
		16'hE6E7: out_word = 8'h66;
		16'hE6E8: out_word = 8'h9D;
		16'hE6E9: out_word = 8'hDE;
		16'hE6EA: out_word = 8'hFB;
		16'hE6EB: out_word = 8'h66;
		16'hE6EC: out_word = 8'hBF;
		16'hE6ED: out_word = 8'h52;
		16'hE6EE: out_word = 8'hB6;
		16'hE6EF: out_word = 8'hFF;
		16'hE6F0: out_word = 8'h66;
		16'hE6F1: out_word = 8'hF5;
		16'hE6F2: out_word = 8'h3E;
		16'hE6F3: out_word = 8'h03;
		16'hE6F4: out_word = 8'hE2;
		16'hE6F5: out_word = 8'hD3;
		16'hE6F6: out_word = 8'h77;
		16'hE6F7: out_word = 8'hAF;
		16'hE6F8: out_word = 8'hD7;
		16'hE6F9: out_word = 8'h57;
		16'hE6FA: out_word = 8'hCC;
		16'hE6FB: out_word = 8'h6D;
		16'hE6FC: out_word = 8'h78;
		16'hE6FD: out_word = 8'h3C;
		16'hE6FE: out_word = 8'h39;
		16'hE6FF: out_word = 8'hAF;
		16'hE700: out_word = 8'hF3;
		16'hE701: out_word = 8'h2F;
		16'hE702: out_word = 8'hF4;
		16'hE703: out_word = 8'hF8;
		16'hE704: out_word = 8'h5B;
		16'hE705: out_word = 8'h09;
		16'hE706: out_word = 8'hEE;
		16'hE707: out_word = 8'h35;
		16'hE708: out_word = 8'hCB;
		16'hE709: out_word = 8'h8D;
		16'hE70A: out_word = 8'hC5;
		16'hE70B: out_word = 8'h6C;
		16'hE70C: out_word = 8'h5F;
		16'hE70D: out_word = 8'hD1;
		16'hE70E: out_word = 8'h5B;
		16'hE70F: out_word = 8'h35;
		16'hE710: out_word = 8'h61;
		16'hE711: out_word = 8'h8D;
		16'hE712: out_word = 8'h7C;
		16'hE713: out_word = 8'h5B;
		16'hE714: out_word = 8'hB4;
		16'hE715: out_word = 8'hE3;
		16'hE716: out_word = 8'h31;
		16'hE717: out_word = 8'hA0;
		16'hE718: out_word = 8'hAF;
		16'hE719: out_word = 8'hD8;
		16'hE71A: out_word = 8'h5B;
		16'hE71B: out_word = 8'h57;
		16'hE71C: out_word = 8'hC7;
		16'hE71D: out_word = 8'hFB;
		16'hE71E: out_word = 8'h5B;
		16'hE71F: out_word = 8'h10;
		16'hE720: out_word = 8'hDB;
		16'hE721: out_word = 8'h57;
		16'hE722: out_word = 8'h18;
		16'hE723: out_word = 8'hFD;
		16'hE724: out_word = 8'h5B;
		16'hE725: out_word = 8'hC5;
		16'hE726: out_word = 8'hCB;
		16'hE727: out_word = 8'hC6;
		16'hE728: out_word = 8'hB2;
		16'hE729: out_word = 8'h8F;
		16'hE72A: out_word = 8'hFD;
		16'hE72B: out_word = 8'hF9;
		16'hE72C: out_word = 8'h6A;
		16'hE72D: out_word = 8'h8B;
		16'hE72E: out_word = 8'h77;
		16'hE72F: out_word = 8'hF0;
		16'hE730: out_word = 8'h80;
		16'hE731: out_word = 8'h61;
		16'hE732: out_word = 8'h8D;
		16'hE733: out_word = 8'h81;
		16'hE734: out_word = 8'h47;
		16'hE735: out_word = 8'h90;
		16'hE736: out_word = 8'hFE;
		16'hE737: out_word = 8'h80;
		16'hE738: out_word = 8'hC5;
		16'hE739: out_word = 8'h0B;
		16'hE73A: out_word = 8'h5F;
		16'hE73B: out_word = 8'hBC;
		16'hE73C: out_word = 8'h80;
		16'hE73D: out_word = 8'h7D;
		16'hE73E: out_word = 8'hBF;
		16'hE73F: out_word = 8'h80;
		16'hE740: out_word = 8'hC3;
		16'hE741: out_word = 8'h14;
		16'hE742: out_word = 8'h25;
		16'hE743: out_word = 8'hF2;
		16'hE744: out_word = 8'h45;
		16'hE745: out_word = 8'hDD;
		16'hE746: out_word = 8'hDC;
		16'hE747: out_word = 8'hDF;
		16'hE748: out_word = 8'hC8;
		16'hE749: out_word = 8'h36;
		16'hE74A: out_word = 8'hE8;
		16'hE74B: out_word = 8'hFE;
		16'hE74C: out_word = 8'h78;
		16'hE74D: out_word = 8'h29;
		16'hE74E: out_word = 8'h8E;
		16'hE74F: out_word = 8'hCB;
		16'hE750: out_word = 8'hFF;
		16'hE751: out_word = 8'h78;
		16'hE752: out_word = 8'h31;
		16'hE753: out_word = 8'h8E;
		16'hE754: out_word = 8'h42;
		16'hE755: out_word = 8'h1A;
		16'hE756: out_word = 8'h75;
		16'hE757: out_word = 8'h24;
		16'hE758: out_word = 8'h77;
		16'hE759: out_word = 8'h2F;
		16'hE75A: out_word = 8'h3E;
		16'hE75B: out_word = 8'hE0;
		16'hE75C: out_word = 8'hE5;
		16'hE75D: out_word = 8'hCD;
		16'hE75E: out_word = 8'h81;
		16'hE75F: out_word = 8'hFA;
		16'hE760: out_word = 8'hE1;
		16'hE761: out_word = 8'hE1;
		16'hE762: out_word = 8'hA7;
		16'hE763: out_word = 8'hCC;
		16'hE764: out_word = 8'h43;
		16'hE765: out_word = 8'hE0;
		16'hE766: out_word = 8'h57;
		16'hE767: out_word = 8'hD5;
		16'hE768: out_word = 8'hF2;
		16'hE769: out_word = 8'h2E;
		16'hE76A: out_word = 8'hFF;
		16'hE76B: out_word = 8'hAF;
		16'hE76C: out_word = 8'h1E;
		16'hE76D: out_word = 8'h1E;
		16'hE76E: out_word = 8'h63;
		16'hE76F: out_word = 8'h7E;
		16'hE770: out_word = 8'hB3;
		16'hE771: out_word = 8'h9D;
		16'hE772: out_word = 8'h26;
		16'hE773: out_word = 8'hFC;
		16'hE774: out_word = 8'h01;
		16'hE775: out_word = 8'h50;
		16'hE776: out_word = 8'hFF;
		16'hE777: out_word = 8'h2E;
		16'hE778: out_word = 8'h0C;
		16'hE779: out_word = 8'h7E;
		16'hE77A: out_word = 8'h87;
		16'hE77B: out_word = 8'h4E;
		16'hE77C: out_word = 8'h06;
		16'hE77D: out_word = 8'hC1;
		16'hE77E: out_word = 8'h0E;
		16'hE77F: out_word = 8'hD0;
		16'hE780: out_word = 8'h40;
		16'hE781: out_word = 8'h04;
		16'hE782: out_word = 8'hB9;
		16'hE783: out_word = 8'hF0;
		16'hE784: out_word = 8'h3E;
		16'hE785: out_word = 8'h91;
		16'hE786: out_word = 8'hFA;
		16'hE787: out_word = 8'hEB;
		16'hE788: out_word = 8'h11;
		16'hE789: out_word = 8'h00;
		16'hE78A: out_word = 8'h10;
		16'hE78B: out_word = 8'h99;
		16'hE78C: out_word = 8'hF8;
		16'hE78D: out_word = 8'h28;
		16'hE78E: out_word = 8'h08;
		16'hE78F: out_word = 8'h69;
		16'hE790: out_word = 8'hF2;
		16'hE791: out_word = 8'hE6;
		16'hE792: out_word = 8'h80;
		16'hE793: out_word = 8'h20;
		16'hE794: out_word = 8'hF5;
		16'hE795: out_word = 8'h34;
		16'hE796: out_word = 8'h53;
		16'hE797: out_word = 8'h2C;
		16'hE798: out_word = 8'hFC;
		16'hE799: out_word = 8'h01;
		16'hE79A: out_word = 8'hC5;
		16'hE79B: out_word = 8'hFA;
		16'hE79C: out_word = 8'hD5;
		16'hE79D: out_word = 8'hCD;
		16'hE79E: out_word = 8'hD6;
		16'hE79F: out_word = 8'h8E;
		16'hE7A0: out_word = 8'h08;
		16'hE7A1: out_word = 8'h5C;
		16'hE7A2: out_word = 8'hDE;
		16'hE7A3: out_word = 8'h20;
		16'hE7A4: out_word = 8'hD8;
		16'hE7A5: out_word = 8'h4A;
		16'hE7A6: out_word = 8'hE4;
		16'hE7A7: out_word = 8'h88;
		16'hE7A8: out_word = 8'h85;
		16'hE7A9: out_word = 8'h4C;
		16'hE7AA: out_word = 8'hF8;
		16'hE7AB: out_word = 8'h37;
		16'hE7AC: out_word = 8'h4F;
		16'hE7AD: out_word = 8'hA6;
		16'hE7AE: out_word = 8'h8E;
		16'hE7AF: out_word = 8'hA5;
		16'hE7B0: out_word = 8'hF1;
		16'hE7B1: out_word = 8'h80;
		16'hE7B2: out_word = 8'h75;
		16'hE7B3: out_word = 8'h3B;
		16'hE7B4: out_word = 8'h4E;
		16'hE7B5: out_word = 8'hF0;
		16'hE7B6: out_word = 8'hD1;
		16'hE7B7: out_word = 8'hC1;
		16'hE7B8: out_word = 8'hB6;
		16'hE7B9: out_word = 8'h9E;
		16'hE7BA: out_word = 8'hB9;
		16'hE7BB: out_word = 8'h2E;
		16'hE7BC: out_word = 8'h40;
		16'hE7BD: out_word = 8'hF8;
		16'hE7BE: out_word = 8'h0E;
		16'hE7BF: out_word = 8'h10;
		16'hE7C0: out_word = 8'hED;
		16'hE7C1: out_word = 8'h58;
		16'hE7C2: out_word = 8'h0C;
		16'hE7C3: out_word = 8'hBF;
		16'hE7C4: out_word = 8'h50;
		16'hE7C5: out_word = 8'h0D;
		16'hE7C6: out_word = 8'h73;
		16'hE7C7: out_word = 8'h23;
		16'hE7C8: out_word = 8'h72;
		16'hE7C9: out_word = 8'h19;
		16'hE7CA: out_word = 8'h8E;
		16'hE7CB: out_word = 8'h0E;
		16'hE7CC: out_word = 8'hF6;
		16'hE7CD: out_word = 8'hC9;
		16'hE7CE: out_word = 8'hD5;
		16'hE7CF: out_word = 8'hC9;
		16'hE7D0: out_word = 8'h37;
		16'hE7D1: out_word = 8'h50;
		16'hE7D2: out_word = 8'h59;
		16'hE7D3: out_word = 8'h01;
		16'hE7D4: out_word = 8'hFB;
		16'hE7D5: out_word = 8'hD0;
		16'hE7D6: out_word = 8'hFF;
		16'hE7D7: out_word = 8'hED;
		16'hE7D8: out_word = 8'h51;
		16'hE7D9: out_word = 8'h08;
		16'hE7DA: out_word = 8'h60;
		16'hE7DB: out_word = 8'hB3;
		16'hE7DC: out_word = 8'h10;
		16'hE7DD: out_word = 8'hB0;
		16'hE7DE: out_word = 8'h30;
		16'hE7DF: out_word = 8'h59;
		16'hE7E0: out_word = 8'hD1;
		16'hE7E1: out_word = 8'hE4;
		16'hE7E2: out_word = 8'h90;
		16'hE7E3: out_word = 8'hEE;
		16'hE7E4: out_word = 8'h49;
		16'hE7E5: out_word = 8'h70;
		16'hE7E6: out_word = 8'hF7;
		16'hE7E7: out_word = 8'h03;
		16'hE7E8: out_word = 8'h50;
		16'hE7E9: out_word = 8'h08;
		16'hE7EA: out_word = 8'h34;
		16'hE7EB: out_word = 8'h8A;
		16'hE7EC: out_word = 8'hC9;
		16'hE7ED: out_word = 8'hDF;
		16'hE7EE: out_word = 8'h68;
		16'hE7EF: out_word = 8'h84;
		16'hE7F0: out_word = 8'hE3;
		16'hE7F1: out_word = 8'hA7;
		16'hE7F2: out_word = 8'h28;
		16'hE7F3: out_word = 8'h3C;
		16'hE7F4: out_word = 8'h8B;
		16'hE7F5: out_word = 8'h39;
		16'hE7F6: out_word = 8'hA5;
		16'hE7F7: out_word = 8'hAF;
		16'hE7F8: out_word = 8'hDD;
		16'hE7F9: out_word = 8'h79;
		16'hE7FA: out_word = 8'h04;
		16'hE7FB: out_word = 8'hDE;
		16'hE7FC: out_word = 8'hCB;
		16'hE7FD: out_word = 8'h3E;
		16'hE7FE: out_word = 8'hEC;
		16'hE7FF: out_word = 8'hEB;
		16'hE800: out_word = 8'h64;
		16'hE801: out_word = 8'hE7;
		16'hE802: out_word = 8'h23;
		16'hE803: out_word = 8'hFC;
		16'hE804: out_word = 8'hE7;
		16'hE805: out_word = 8'h20;
		16'hE806: out_word = 8'h3D;
		16'hE807: out_word = 8'h0F;
		16'hE808: out_word = 8'h38;
		16'hE809: out_word = 8'h07;
		16'hE80A: out_word = 8'h77;
		16'hE80B: out_word = 8'hA9;
		16'hE80C: out_word = 8'h60;
		16'hE80D: out_word = 8'hED;
		16'hE80E: out_word = 8'hE1;
		16'hE80F: out_word = 8'h58;
		16'hE810: out_word = 8'h49;
		16'hE811: out_word = 8'hD9;
		16'hE812: out_word = 8'h50;
		16'hE813: out_word = 8'h30;
		16'hE814: out_word = 8'h9D;
		16'hE815: out_word = 8'hCA;
		16'hE816: out_word = 8'h58;
		16'hE817: out_word = 8'h21;
		16'hE818: out_word = 8'h14;
		16'hE819: out_word = 8'h4C;
		16'hE81A: out_word = 8'h34;
		16'hE81B: out_word = 8'hCB;
		16'hE81C: out_word = 8'h36;
		16'hE81D: out_word = 8'hC8;
		16'hE81E: out_word = 8'h2F;
		16'hE81F: out_word = 8'h7F;
		16'hE820: out_word = 8'h6C;
		16'hE821: out_word = 8'h45;
		16'hE822: out_word = 8'h5C;
		16'hE823: out_word = 8'h8F;
		16'hE824: out_word = 8'hBF;
		16'hE825: out_word = 8'hF1;
		16'hE826: out_word = 8'hCD;
		16'hE827: out_word = 8'h64;
		16'hE828: out_word = 8'h8F;
		16'hE829: out_word = 8'hA7;
		16'hE82A: out_word = 8'hA2;
		16'hE82B: out_word = 8'hDE;
		16'hE82C: out_word = 8'h42;
		16'hE82D: out_word = 8'hE0;
		16'hE82E: out_word = 8'hFF;
		16'hE82F: out_word = 8'hE5;
		16'hE830: out_word = 8'hEB;
		16'hE831: out_word = 8'h21;
		16'hE832: out_word = 8'hF0;
		16'hE833: out_word = 8'h3F;
		16'hE834: out_word = 8'h01;
		16'hE835: out_word = 8'h06;
		16'hE836: out_word = 8'h00;
		16'hE837: out_word = 8'hF0;
		16'hE838: out_word = 8'hCD;
		16'hE839: out_word = 8'h76;
		16'hE83A: out_word = 8'h90;
		16'hE83B: out_word = 8'hE1;
		16'hE83C: out_word = 8'h81;
		16'hE83D: out_word = 8'hC2;
		16'hE83E: out_word = 8'h11;
		16'hE83F: out_word = 8'h7E;
		16'hE840: out_word = 8'hF9;
		16'hE841: out_word = 8'h1A;
		16'hE842: out_word = 8'hBE;
		16'hE843: out_word = 8'h13;
		16'hE844: out_word = 8'h23;
		16'hE845: out_word = 8'h20;
		16'hE846: out_word = 8'h2E;
		16'hE847: out_word = 8'hF8;
		16'hE848: out_word = 8'hF8;
		16'hE849: out_word = 8'h01;
		16'hE84A: out_word = 8'hBA;
		16'hE84B: out_word = 8'h5F;
		16'hE84C: out_word = 8'h3B;
		16'hE84D: out_word = 8'hFF;
		16'hE84E: out_word = 8'hE1;
		16'hE84F: out_word = 8'hCD;
		16'hE850: out_word = 8'h84;
		16'hE851: out_word = 8'h90;
		16'hE852: out_word = 8'h3C;
		16'hE853: out_word = 8'hF5;
		16'hE854: out_word = 8'h20;
		16'hE855: out_word = 8'h05;
		16'hE856: out_word = 8'h21;
		16'hE857: out_word = 8'hFF;
		16'hE858: out_word = 8'hF2;
		16'hE859: out_word = 8'hB5;
		16'hE85A: out_word = 8'hEF;
		16'hE85B: out_word = 8'h12;
		16'hE85C: out_word = 8'hF7;
		16'hE85D: out_word = 8'h56;
		16'hE85E: out_word = 8'h6E;
		16'hE85F: out_word = 8'h90;
		16'hE860: out_word = 8'hE5;
		16'hE861: out_word = 8'h0A;
		16'hE862: out_word = 8'hE0;
		16'hE863: out_word = 8'h14;
		16'hE864: out_word = 8'h8C;
		16'hE865: out_word = 8'h25;
		16'hE866: out_word = 8'hFD;
		16'hE867: out_word = 8'h9B;
		16'hE868: out_word = 8'hA8;
		16'hE869: out_word = 8'h8F;
		16'hE86A: out_word = 8'h99;
		16'hE86B: out_word = 8'hFF;
		16'hE86C: out_word = 8'h9B;
		16'hE86D: out_word = 8'h2A;
		16'hE86E: out_word = 8'h01;
		16'hE86F: out_word = 8'hBE;
		16'hE870: out_word = 8'hFA;
		16'hE871: out_word = 8'h5F;
		16'hE872: out_word = 8'h9B;
		16'hE873: out_word = 8'h40;
		16'hE874: out_word = 8'hDD;
		16'hE875: out_word = 8'h8C;
		16'hE876: out_word = 8'hB6;
		16'hE877: out_word = 8'hFE;
		16'hE878: out_word = 8'h0A;
		16'hE879: out_word = 8'h3D;
		16'hE87A: out_word = 8'h00;
		16'hE87B: out_word = 8'hF7;
		16'hE87C: out_word = 8'h68;
		16'hE87D: out_word = 8'hCD;
		16'hE87E: out_word = 8'h91;
		16'hE87F: out_word = 8'hF9;
		16'hE880: out_word = 8'hD7;
		16'hE881: out_word = 8'hF4;
		16'hE882: out_word = 8'h98;
		16'hE883: out_word = 8'h09;
		16'hE884: out_word = 8'hB2;
		16'hE885: out_word = 8'h4B;
		16'hE886: out_word = 8'h0F;
		16'hE887: out_word = 8'hF4;
		16'hE888: out_word = 8'h27;
		16'hE889: out_word = 8'hFD;
		16'hE88A: out_word = 8'h97;
		16'hE88B: out_word = 8'h4D;
		16'hE88C: out_word = 8'h90;
		16'hE88D: out_word = 8'h08;
		16'hE88E: out_word = 8'h2F;
		16'hE88F: out_word = 8'hDC;
		16'hE890: out_word = 8'h20;
		16'hE891: out_word = 8'h23;
		16'hE892: out_word = 8'hD5;
		16'hE893: out_word = 8'hE2;
		16'hE894: out_word = 8'hD1;
		16'hE895: out_word = 8'h35;
		16'hE896: out_word = 8'hF7;
		16'hE897: out_word = 8'h7B;
		16'hE898: out_word = 8'hF5;
		16'hE899: out_word = 8'hCD;
		16'hE89A: out_word = 8'h12;
		16'hE89B: out_word = 8'h51;
		16'hE89C: out_word = 8'hF0;
		16'hE89D: out_word = 8'hD2;
		16'hE89E: out_word = 8'hD7;
		16'hE89F: out_word = 8'hF9;
		16'hE8A0: out_word = 8'hF1;
		16'hE8A1: out_word = 8'h5B;
		16'hE8A2: out_word = 8'hC0;
		16'hE8A3: out_word = 8'h7F;
		16'hE8A4: out_word = 8'h94;
		16'hE8A5: out_word = 8'h11;
		16'hE8A6: out_word = 8'hD8;
		16'hE8A7: out_word = 8'hFA;
		16'hE8A8: out_word = 8'hF8;
		16'hE8A9: out_word = 8'h3E;
		16'hE8AA: out_word = 8'h40;
		16'hE8AB: out_word = 8'h08;
		16'hE8AC: out_word = 8'h42;
		16'hE8AD: out_word = 8'h77;
		16'hE8AE: out_word = 8'hE6;
		16'hE8AF: out_word = 8'h77;
		16'hE8B0: out_word = 8'h23;
		16'hE8B1: out_word = 8'h43;
		16'hE8B2: out_word = 8'h98;
		16'hE8B3: out_word = 8'hFA;
		16'hE8B4: out_word = 8'h44;
		16'hE8B5: out_word = 8'hF4;
		16'hE8B6: out_word = 8'h5F;
		16'hE8B7: out_word = 8'h52;
		16'hE8B8: out_word = 8'hBB;
		16'hE8B9: out_word = 8'hCB;
		16'hE8BA: out_word = 8'hE0;
		16'hE8BB: out_word = 8'h89;
		16'hE8BC: out_word = 8'h1D;
		16'hE8BD: out_word = 8'h5F;
		16'hE8BE: out_word = 8'hFE;
		16'hE8BF: out_word = 8'h7A;
		16'hE8C0: out_word = 8'hCD;
		16'hE8C1: out_word = 8'h95;
		16'hE8C2: out_word = 8'hFD;
		16'hE8C3: out_word = 8'h7B;
		16'hE8C4: out_word = 8'h20;
		16'hE8C5: out_word = 8'hFA;
		16'hE8C6: out_word = 8'hD1;
		16'hE8C7: out_word = 8'hDE;
		16'hE8C8: out_word = 8'hFC;
		16'hE8C9: out_word = 8'hF3;
		16'hE8CA: out_word = 8'hB8;
		16'hE8CB: out_word = 8'hFB;
		16'hE8CC: out_word = 8'hF3;
		16'hE8CD: out_word = 8'h17;
		16'hE8CE: out_word = 8'hFA;
		16'hE8CF: out_word = 8'h08;
		16'hE8D0: out_word = 8'hE5;
		16'hE8D1: out_word = 8'h5F;
		16'hE8D2: out_word = 8'hF7;
		16'hE8D3: out_word = 8'hAB;
		16'hE8D4: out_word = 8'hE3;
		16'hE8D5: out_word = 8'h1D;
		16'hE8D6: out_word = 8'hEB;
		16'hE8D7: out_word = 8'hF8;
		16'hE8D8: out_word = 8'h0D;
		16'hE8D9: out_word = 8'h18;
		16'hE8DA: out_word = 8'hC5;
		16'hE8DB: out_word = 8'hF8;
		16'hE8DC: out_word = 8'hF5;
		16'hE8DD: out_word = 8'h79;
		16'hE8DE: out_word = 8'hC3;
		16'hE8DF: out_word = 8'hBB;
		16'hE8E0: out_word = 8'hF2;
		16'hE8E1: out_word = 8'hF3;
		16'hE8E2: out_word = 8'h79;
		16'hE8E3: out_word = 8'hEA;
		16'hE8E4: out_word = 8'h1E;
		16'hE8E5: out_word = 8'hC5;
		16'hE8E6: out_word = 8'h5B;
		16'hE8E7: out_word = 8'hD6;
		16'hE8E8: out_word = 8'h16;
		16'hE8E9: out_word = 8'h1A;
		16'hE8EA: out_word = 8'hBA;
		16'hE8EB: out_word = 8'h90;
		16'hE8EC: out_word = 8'h15;
		16'hE8ED: out_word = 8'h28;
		16'hE8EE: out_word = 8'h4D;
		16'hE8EF: out_word = 8'h7F;
		16'hE8F0: out_word = 8'hA7;
		16'hE8F1: out_word = 8'hCB;
		16'hE8F2: out_word = 8'h7F;
		16'hE8F3: out_word = 8'h20;
		16'hE8F4: out_word = 8'hF3;
		16'hE8F5: out_word = 8'hA7;
		16'hE8F6: out_word = 8'h28;
		16'hE8F7: out_word = 8'h43;
		16'hE8F8: out_word = 8'h8B;
		16'hE8F9: out_word = 8'h3C;
		16'hE8FA: out_word = 8'h40;
		16'hE8FB: out_word = 8'h94;
		16'hE8FC: out_word = 8'hAF;
		16'hE8FD: out_word = 8'hAE;
		16'hE8FE: out_word = 8'hE3;
		16'hE8FF: out_word = 8'h29;
		16'hE900: out_word = 8'hB0;
		16'hE901: out_word = 8'hFB;
		16'hE902: out_word = 8'h3E;
		16'hE903: out_word = 8'h96;
		16'hE904: out_word = 8'hEC;
		16'hE905: out_word = 8'hDC;
		16'hE906: out_word = 8'hC3;
		16'hE907: out_word = 8'h32;
		16'hE908: out_word = 8'hE3;
		16'hE909: out_word = 8'h26;
		16'hE90A: out_word = 8'h36;
		16'hE90B: out_word = 8'hE3;
		16'hE90C: out_word = 8'h23;
		16'hE90D: out_word = 8'h47;
		16'hE90E: out_word = 8'hE5;
		16'hE90F: out_word = 8'h5C;
		16'hE910: out_word = 8'hEC;
		16'hE911: out_word = 8'hDE;
		16'hE912: out_word = 8'h25;
		16'hE913: out_word = 8'hEA;
		16'hE914: out_word = 8'h5F;
		16'hE915: out_word = 8'hD3;
		16'hE916: out_word = 8'h39;
		16'hE917: out_word = 8'hFA;
		16'hE918: out_word = 8'h57;
		16'hE919: out_word = 8'hB3;
		16'hE91A: out_word = 8'hCA;
		16'hE91B: out_word = 8'h1C;
		16'hE91C: out_word = 8'h5F;
		16'hE91D: out_word = 8'h59;
		16'hE91E: out_word = 8'hF5;
		16'hE91F: out_word = 8'h3E;
		16'hE920: out_word = 8'h01;
		16'hE921: out_word = 8'hED;
		16'hE922: out_word = 8'h52;
		16'hE923: out_word = 8'hF6;
		16'hE924: out_word = 8'h59;
		16'hE925: out_word = 8'h4D;
		16'hE926: out_word = 8'hFC;
		16'hE927: out_word = 8'h23;
		16'hE928: out_word = 8'hED;
		16'hE929: out_word = 8'h73;
		16'hE92A: out_word = 8'h00;
		16'hE92B: out_word = 8'hD7;
		16'hE92C: out_word = 8'h13;
		16'hE92D: out_word = 8'hE6;
		16'hE92E: out_word = 8'h91;
		16'hE92F: out_word = 8'h57;
		16'hE930: out_word = 8'h1F;
		16'hE931: out_word = 8'h86;
		16'hE932: out_word = 8'h19;
		16'hE933: out_word = 8'hCB;
		16'hE934: out_word = 8'hFE;
		16'hE935: out_word = 8'h4C;
		16'hE936: out_word = 8'hED;
		16'hE937: out_word = 8'h7B;
		16'hE938: out_word = 8'h5F;
		16'hE939: out_word = 8'hE6;
		16'hE93A: out_word = 8'h7F;
		16'hE93B: out_word = 8'h1B;
		16'hE93C: out_word = 8'hA4;
		16'hE93D: out_word = 8'h94;
		16'hE93E: out_word = 8'hBC;
		16'hE93F: out_word = 8'h92;
		16'hE940: out_word = 8'h8D;
		16'hE941: out_word = 8'h56;
		16'hE942: out_word = 8'hC5;
		16'hE943: out_word = 8'hC6;
		16'hE944: out_word = 8'h91;
		16'hE945: out_word = 8'h2D;
		16'hE946: out_word = 8'hFE;
		16'hE947: out_word = 8'h1E;
		16'hE948: out_word = 8'h96;
		16'hE949: out_word = 8'h7C;
		16'hE94A: out_word = 8'h93;
		16'hE94B: out_word = 8'h71;
		16'hE94C: out_word = 8'h94;
		16'hE94D: out_word = 8'h52;
		16'hE94E: out_word = 8'h37;
		16'hE94F: out_word = 8'h0B;
		16'hE950: out_word = 8'h98;
		16'hE951: out_word = 8'hD9;
		16'hE952: out_word = 8'hC5;
		16'hE953: out_word = 8'h1E;
		16'hE954: out_word = 8'h00;
		16'hE955: out_word = 8'hFF;
		16'hE956: out_word = 8'hF5;
		16'hE957: out_word = 8'hE5;
		16'hE958: out_word = 8'h08;
		16'hE959: out_word = 8'h3A;
		16'hE95A: out_word = 8'h04;
		16'hE95B: out_word = 8'hD7;
		16'hE95C: out_word = 8'h67;
		16'hE95D: out_word = 8'hD5;
		16'hE95E: out_word = 8'hFF;
		16'hE95F: out_word = 8'hCD;
		16'hE960: out_word = 8'hAA;
		16'hE961: out_word = 8'h97;
		16'hE962: out_word = 8'h4C;
		16'hE963: out_word = 8'h21;
		16'hE964: out_word = 8'h00;
		16'hE965: out_word = 8'hD8;
		16'hE966: out_word = 8'hEB;
		16'hE967: out_word = 8'h56;
		16'hE968: out_word = 8'h28;
		16'hE969: out_word = 8'h13;
		16'hE96A: out_word = 8'hE1;
		16'hE96B: out_word = 8'h79;
		16'hE96C: out_word = 8'hFE;
		16'hE96D: out_word = 8'h06;
		16'hE96E: out_word = 8'h00;
		16'hE96F: out_word = 8'h3D;
		16'hE970: out_word = 8'hA5;
		16'hE971: out_word = 8'h28;
		16'hE972: out_word = 8'h19;
		16'hE973: out_word = 8'hD9;
		16'hE974: out_word = 8'hA0;
		16'hE975: out_word = 8'hFC;
		16'hE976: out_word = 8'h27;
		16'hE977: out_word = 8'h6F;
		16'hE978: out_word = 8'h79;
		16'hE979: out_word = 8'h95;
		16'hE97A: out_word = 8'hFF;
		16'hE97B: out_word = 8'h67;
		16'hE97C: out_word = 8'h08;
		16'hE97D: out_word = 8'hBC;
		16'hE97E: out_word = 8'h38;
		16'hE97F: out_word = 8'h01;
		16'hE980: out_word = 8'h7C;
		16'hE981: out_word = 8'hE1;
		16'hE982: out_word = 8'hE5;
		16'hE983: out_word = 8'hF4;
		16'hE984: out_word = 8'hCD;
		16'hE985: out_word = 8'hBE;
		16'hE986: out_word = 8'h91;
		16'hE987: out_word = 8'h41;
		16'hE988: out_word = 8'hD3;
		16'hE989: out_word = 8'hF9;
		16'hE98A: out_word = 8'h4F;
		16'hE98B: out_word = 8'hE3;
		16'hE98C: out_word = 8'hD9;
		16'hE98D: out_word = 8'h01;
		16'hE98E: out_word = 8'h00;
		16'hE98F: out_word = 8'hE7;
		16'hE990: out_word = 8'hF3;
		16'hE991: out_word = 8'hE1;
		16'hE992: out_word = 8'hF1;
		16'hE993: out_word = 8'h90;
		16'hE994: out_word = 8'hC8;
		16'hE995: out_word = 8'hE0;
		16'hE996: out_word = 8'hB9;
		16'hE997: out_word = 8'hFF;
		16'hE998: out_word = 8'h28;
		16'hE999: out_word = 8'h4A;
		16'hE99A: out_word = 8'h04;
		16'hE99B: out_word = 8'h91;
		16'hE99C: out_word = 8'h30;
		16'hE99D: out_word = 8'hFC;
		16'hE99E: out_word = 8'h05;
		16'hE99F: out_word = 8'h81;
		16'hE9A0: out_word = 8'hAF;
		16'hE9A1: out_word = 8'hF5;
		16'hE9A2: out_word = 8'h61;
		16'hE9A3: out_word = 8'hA0;
		16'hE9A4: out_word = 8'h3E;
		16'hE9A5: out_word = 8'hF1;
		16'hE9A6: out_word = 8'h7F;
		16'hE9A7: out_word = 8'hC5;
		16'hE9A8: out_word = 8'hE5;
		16'hE9A9: out_word = 8'h79;
		16'hE9AA: out_word = 8'hEB;
		16'hE9AB: out_word = 8'hCD;
		16'hE9AC: out_word = 8'h9B;
		16'hE9AD: out_word = 8'h94;
		16'hE9AE: out_word = 8'hF4;
		16'hE9AF: out_word = 8'hCB;
		16'hE9B0: out_word = 8'h78;
		16'hE9B1: out_word = 8'hC2;
		16'hE9B2: out_word = 8'h10;
		16'hE9B3: out_word = 8'h71;
		16'hE9B4: out_word = 8'hFC;
		16'hE9B5: out_word = 8'hF5;
		16'hE9B6: out_word = 8'hCD;
		16'hE9B7: out_word = 8'h59;
		16'hE9B8: out_word = 8'h97;
		16'hE9B9: out_word = 8'hD9;
		16'hE9BA: out_word = 8'hC5;
		16'hE9BB: out_word = 8'h95;
		16'hE9BC: out_word = 8'hD5;
		16'hE9BD: out_word = 8'hAC;
		16'hE9BE: out_word = 8'hCF;
		16'hE9BF: out_word = 8'h45;
		16'hE9C0: out_word = 8'hED;
		16'hE9C1: out_word = 8'h4A;
		16'hE9C2: out_word = 8'h44;
		16'hE9C3: out_word = 8'h4D;
		16'hE9C4: out_word = 8'hF8;
		16'hE9C5: out_word = 8'hF1;
		16'hE9C6: out_word = 8'hE1;
		16'hE9C7: out_word = 8'h08;
		16'hE9C8: out_word = 8'hD9;
		16'hE9C9: out_word = 8'h7B;
		16'hE9CA: out_word = 8'hC6;
		16'hE9CB: out_word = 8'hD6;
		16'hE9CC: out_word = 8'h07;
		16'hE9CD: out_word = 8'h0F;
		16'hE9CE: out_word = 8'hCD;
		16'hE9CF: out_word = 8'h09;
		16'hE9D0: out_word = 8'h87;
		16'hE9D1: out_word = 8'hC6;
		16'hE9D2: out_word = 8'h05;
		16'hE9D3: out_word = 8'h18;
		16'hE9D4: out_word = 8'h73;
		16'hE9D5: out_word = 8'hF9;
		16'hE9D6: out_word = 8'h03;
		16'hE9D7: out_word = 8'hA7;
		16'hE9D8: out_word = 8'h4C;
		16'hE9D9: out_word = 8'hD4;
		16'hE9DA: out_word = 8'hD1;
		16'hE9DB: out_word = 8'hC1;
		16'hE9DC: out_word = 8'h4F;
		16'hE9DD: out_word = 8'hC4;
		16'hE9DE: out_word = 8'hF1;
		16'hE9DF: out_word = 8'h04;
		16'hE9E0: out_word = 8'hA7;
		16'hE9E1: out_word = 8'hFC;
		16'hE9E2: out_word = 8'hC8;
		16'hE9E3: out_word = 8'h4F;
		16'hE9E4: out_word = 8'hAF;
		16'hE9E5: out_word = 8'h18;
		16'hE9E6: out_word = 8'hBB;
		16'hE9E7: out_word = 8'hCD;
		16'hE9E8: out_word = 8'hFA;
		16'hE9E9: out_word = 8'h55;
		16'hE9EA: out_word = 8'h11;
		16'hE9EB: out_word = 8'h14;
		16'hE9EC: out_word = 8'h00;
		16'hE9ED: out_word = 8'h19;
		16'hE9EE: out_word = 8'hA6;
		16'hE9EF: out_word = 8'h05;
		16'hE9F0: out_word = 8'h1E;
		16'hE9F1: out_word = 8'h05;
		16'hE9F2: out_word = 8'hED;
		16'hE9F3: out_word = 8'h00;
		16'hE9F4: out_word = 8'h05;
		16'hE9F5: out_word = 8'hBE;
		16'hE9F6: out_word = 8'h0A;
		16'hE9F7: out_word = 8'h7C;
		16'hE9F8: out_word = 8'hAD;
		16'hE9F9: out_word = 8'hED;
		16'hE9FA: out_word = 8'h53;
		16'hE9FB: out_word = 8'h25;
		16'hE9FC: out_word = 8'hD7;
		16'hE9FD: out_word = 8'h4C;
		16'hE9FE: out_word = 8'h43;
		16'hE9FF: out_word = 8'h27;
		16'hEA00: out_word = 8'h42;
		16'hEA01: out_word = 8'hD6;
		16'hEA02: out_word = 8'h9C;
		16'hEA03: out_word = 8'h58;
		16'hEA04: out_word = 8'hCD;
		16'hEA05: out_word = 8'h92;
		16'hEA06: out_word = 8'h94;
		16'hEA07: out_word = 8'h87;
		16'hEA08: out_word = 8'h71;
		16'hEA09: out_word = 8'h96;
		16'hEA0A: out_word = 8'h06;
		16'hEA0B: out_word = 8'hAC;
		16'hEA0C: out_word = 8'h2F;
		16'hEA0D: out_word = 8'hE1;
		16'hEA0E: out_word = 8'h30;
		16'hEA0F: out_word = 8'hF3;
		16'hEA10: out_word = 8'h5F;
		16'hEA11: out_word = 8'hC6;
		16'hEA12: out_word = 8'h9A;
		16'hEA13: out_word = 8'h92;
		16'hEA14: out_word = 8'hE1;
		16'hEA15: out_word = 8'h5B;
		16'hEA16: out_word = 8'h4F;
		16'hEA17: out_word = 8'hE1;
		16'hEA18: out_word = 8'h4B;
		16'hEA19: out_word = 8'hE1;
		16'hEA1A: out_word = 8'hCD;
		16'hEA1B: out_word = 8'h08;
		16'hEA1C: out_word = 8'h92;
		16'hEA1D: out_word = 8'hFF;
		16'hEA1E: out_word = 8'hC3;
		16'hEA1F: out_word = 8'h99;
		16'hEA20: out_word = 8'h97;
		16'hEA21: out_word = 8'h7A;
		16'hEA22: out_word = 8'hE6;
		16'hEA23: out_word = 8'h01;
		16'hEA24: out_word = 8'h67;
		16'hEA25: out_word = 8'h7B;
		16'hEA26: out_word = 8'h21;
		16'hEA27: out_word = 8'h99;
		16'hEA28: out_word = 8'hCF;
		16'hEA29: out_word = 8'h24;
		16'hEA2A: out_word = 8'h1D;
		16'hEA2B: out_word = 8'h6B;
		16'hEA2C: out_word = 8'hCB;
		16'hEA2D: out_word = 8'h44;
		16'hEA2E: out_word = 8'h40;
		16'hEA2F: out_word = 8'hF8;
		16'hEA30: out_word = 8'hED;
		16'hEA31: out_word = 8'h82;
		16'hEA32: out_word = 8'hD8;
		16'hEA33: out_word = 8'h7C;
		16'hEA34: out_word = 8'hC9;
		16'hEA35: out_word = 8'hCD;
		16'hEA36: out_word = 8'h9D;
		16'hEA37: out_word = 8'h92;
		16'hEA38: out_word = 8'h20;
		16'hEA39: out_word = 8'h04;
		16'hEA3A: out_word = 8'h5A;
		16'hEA3B: out_word = 8'h87;
		16'hEA3C: out_word = 8'hC9;
		16'hEA3D: out_word = 8'h73;
		16'hEA3E: out_word = 8'hB1;
		16'hEA3F: out_word = 8'h33;
		16'hEA40: out_word = 8'hD7;
		16'hEA41: out_word = 8'hA9;
		16'hEA42: out_word = 8'h31;
		16'hEA43: out_word = 8'h11;
		16'hEA44: out_word = 8'h29;
		16'hEA45: out_word = 8'hF4;
		16'hEA46: out_word = 8'hE5;
		16'hEA47: out_word = 8'h77;
		16'hEA48: out_word = 8'h02;
		16'hEA49: out_word = 8'h73;
		16'hEA4A: out_word = 8'h77;
		16'hEA4B: out_word = 8'hE1;
		16'hEA4C: out_word = 8'hC9;
		16'hEA4D: out_word = 8'h9F;
		16'hEA4E: out_word = 8'h21;
		16'hEA4F: out_word = 8'hEF;
		16'hEA50: out_word = 8'h7E;
		16'hEA51: out_word = 8'h23;
		16'hEA52: out_word = 8'hBB;
		16'hEA53: out_word = 8'hC0;
		16'hEA54: out_word = 8'h34;
		16'hEA55: out_word = 8'hFC;
		16'hEA56: out_word = 8'hBA;
		16'hEA57: out_word = 8'hFC;
		16'hEA58: out_word = 8'h9D;
		16'hEA59: out_word = 8'hB9;
		16'hEA5A: out_word = 8'hFC;
		16'hEA5B: out_word = 8'hB8;
		16'hEA5C: out_word = 8'hC9;
		16'hEA5D: out_word = 8'h3C;
		16'hEA5E: out_word = 8'h6F;
		16'hEA5F: out_word = 8'hCB;
		16'hEA60: out_word = 8'h67;
		16'hEA61: out_word = 8'h08;
		16'hEA62: out_word = 8'h7B;
		16'hEA63: out_word = 8'h6F;
		16'hEA64: out_word = 8'h5F;
		16'hEA65: out_word = 8'h56;
		16'hEA66: out_word = 8'hC8;
		16'hEA67: out_word = 8'hD9;
		16'hEA68: out_word = 8'h07;
		16'hEA69: out_word = 8'hCB;
		16'hEA6A: out_word = 8'h7F;
		16'hEA6B: out_word = 8'hF3;
		16'hEA6C: out_word = 8'h28;
		16'hEA6D: out_word = 8'h14;
		16'hEA6E: out_word = 8'h21;
		16'hEA6F: out_word = 8'h3E;
		16'hEA70: out_word = 8'hDD;
		16'hEA71: out_word = 8'hA7;
		16'hEA72: out_word = 8'h9F;
		16'hEA73: out_word = 8'hD9;
		16'hEA74: out_word = 8'hF3;
		16'hEA75: out_word = 8'h3D;
		16'hEA76: out_word = 8'h77;
		16'hEA77: out_word = 8'h87;
		16'hEA78: out_word = 8'h26;
		16'hEA79: out_word = 8'hF8;
		16'hEA7A: out_word = 8'hD6;
		16'hEA7B: out_word = 8'h6F;
		16'hEA7C: out_word = 8'h7E;
		16'hEA7D: out_word = 8'h2C;
		16'hEA7E: out_word = 8'h66;
		16'hEA7F: out_word = 8'h9B;
		16'hEA80: out_word = 8'h18;
		16'hEA81: out_word = 8'h17;
		16'hEA82: out_word = 8'h9D;
		16'hEA83: out_word = 8'hEC;
		16'hEA84: out_word = 8'h3C;
		16'hEA85: out_word = 8'hFE;
		16'hEA86: out_word = 8'h80;
		16'hEA87: out_word = 8'h37;
		16'hEA88: out_word = 8'hEA;
		16'hEA89: out_word = 8'h77;
		16'hEA8A: out_word = 8'h3D;
		16'hEA8B: out_word = 8'h0F;
		16'hEA8C: out_word = 8'hEA;
		16'hEA8D: out_word = 8'h73;
		16'hEA8E: out_word = 8'h39;
		16'hEA8F: out_word = 8'hD7;
		16'hEA90: out_word = 8'h71;
		16'hEA91: out_word = 8'hF6;
		16'hEA92: out_word = 8'h2C;
		16'hEA93: out_word = 8'h70;
		16'hEA94: out_word = 8'hD9;
		16'hEA95: out_word = 8'hD5;
		16'hEA96: out_word = 8'h5B;
		16'hEA97: out_word = 8'h34;
		16'hEA98: out_word = 8'h78;
		16'hEA99: out_word = 8'hB1;
		16'hEA9A: out_word = 8'hF3;
		16'hEA9B: out_word = 8'hB2;
		16'hEA9C: out_word = 8'hB3;
		16'hEA9D: out_word = 8'h20;
		16'hEA9E: out_word = 8'h08;
		16'hEA9F: out_word = 8'h53;
		16'hEAA0: out_word = 8'h05;
		16'hEAA1: out_word = 8'h4A;
		16'hEAA2: out_word = 8'h53;
		16'hEAA3: out_word = 8'h07;
		16'hEAA4: out_word = 8'h52;
		16'hEAA5: out_word = 8'h83;
		16'hEAA6: out_word = 8'h35;
		16'hEAA7: out_word = 8'h2C;
		16'hEAA8: out_word = 8'h37;
		16'hEAA9: out_word = 8'h7D;
		16'hEAAA: out_word = 8'h4B;
		16'hEAAB: out_word = 8'h3D;
		16'hEAAC: out_word = 8'h93;
		16'hEAAD: out_word = 8'hD1;
		16'hEAAE: out_word = 8'hC9;
		16'hEAAF: out_word = 8'hC3;
		16'hEAB0: out_word = 8'hCF;
		16'hEAB1: out_word = 8'hE1;
		16'hEAB2: out_word = 8'h28;
		16'hEAB3: out_word = 8'hFF;
		16'hEAB4: out_word = 8'h07;
		16'hEAB5: out_word = 8'hC5;
		16'hEAB6: out_word = 8'h0B;
		16'hEAB7: out_word = 8'hCD;
		16'hEAB8: out_word = 8'hCB;
		16'hEAB9: out_word = 8'h92;
		16'hEABA: out_word = 8'hC1;
		16'hEABB: out_word = 8'h5F;
		16'hEABC: out_word = 8'h30;
		16'hEABD: out_word = 8'h0C;
		16'hEABE: out_word = 8'hFB;
		16'hEABF: out_word = 8'hBF;
		16'hEAC0: out_word = 8'hD1;
		16'hEAC1: out_word = 8'h3C;
		16'hEAC2: out_word = 8'h7B;
		16'hEAC3: out_word = 8'hC8;
		16'hEAC4: out_word = 8'h08;
		16'hEAC5: out_word = 8'h79;
		16'hEAC6: out_word = 8'hD6;
		16'hEAC7: out_word = 8'hE6;
		16'hEAC8: out_word = 8'h0F;
		16'hEAC9: out_word = 8'h17;
		16'hEACA: out_word = 8'hF9;
		16'hEACB: out_word = 8'hDF;
		16'hEACC: out_word = 8'h66;
		16'hEACD: out_word = 8'h3F;
		16'hEACE: out_word = 8'h41;
		16'hEACF: out_word = 8'h0B;
		16'hEAD0: out_word = 8'h00;
		16'hEAD1: out_word = 8'h7E;
		16'hEAD2: out_word = 8'hEB;
		16'hEAD3: out_word = 8'h0B;
		16'hEAD4: out_word = 8'h6E;
		16'hEAD5: out_word = 8'h67;
		16'hEAD6: out_word = 8'h13;
		16'hEAD7: out_word = 8'hCD;
		16'hEAD8: out_word = 8'h70;
		16'hEAD9: out_word = 8'hD4;
		16'hEADA: out_word = 8'h93;
		16'hEADB: out_word = 8'h16;
		16'hEADC: out_word = 8'h84;
		16'hEADD: out_word = 8'hFF;
		16'hEADE: out_word = 8'hFF;
		16'hEADF: out_word = 8'h80;
		16'hEAE0: out_word = 8'h08;
		16'hEAE1: out_word = 8'hFE;
		16'hEAE2: out_word = 8'h0F;
		16'hEAE3: out_word = 8'h7B;
		16'hEAE4: out_word = 8'h5A;
		16'hEAE5: out_word = 8'hC0;
		16'hEAE6: out_word = 8'h1C;
		16'hEAE7: out_word = 8'hD7;
		16'hEAE8: out_word = 8'hC9;
		16'hEAE9: out_word = 8'hC5;
		16'hEAEA: out_word = 8'h0E;
		16'hEAEB: out_word = 8'hDB;
		16'hEAEC: out_word = 8'h1F;
		16'hEAED: out_word = 8'h3E;
		16'hEAEE: out_word = 8'h10;
		16'hEAEF: out_word = 8'hBF;
		16'hEAF0: out_word = 8'h36;
		16'hEAF1: out_word = 8'h7B;
		16'hEAF2: out_word = 8'hAF;
		16'hEAF3: out_word = 8'hF5;
		16'hEAF4: out_word = 8'h88;
		16'hEAF5: out_word = 8'h59;
		16'hEAF6: out_word = 8'h86;
		16'hEAF7: out_word = 8'hF7;
		16'hEAF8: out_word = 8'h27;
		16'hEAF9: out_word = 8'hD2;
		16'hEAFA: out_word = 8'hEF;
		16'hEAFB: out_word = 8'hBF;
		16'hEAFC: out_word = 8'h2E;
		16'hEAFD: out_word = 8'hFC;
		16'hEAFE: out_word = 8'h6F;
		16'hEAFF: out_word = 8'h28;
		16'hEB00: out_word = 8'h06;
		16'hEB01: out_word = 8'hC1;
		16'hEB02: out_word = 8'hF5;
		16'hEB03: out_word = 8'hFF;
		16'hEB04: out_word = 8'hAF;
		16'hEB05: out_word = 8'h3D;
		16'hEB06: out_word = 8'hC9;
		16'hEB07: out_word = 8'hF8;
		16'hEB08: out_word = 8'h6D;
		16'hEB09: out_word = 8'hF1;
		16'hEB0A: out_word = 8'h51;
		16'hEB0B: out_word = 8'h6F;
		16'hEB0C: out_word = 8'h6A;
		16'hEB0D: out_word = 8'hA5;
		16'hEB0E: out_word = 8'hCD;
		16'hEB0F: out_word = 8'hCA;
		16'hEB10: out_word = 8'hFF;
		16'hEB11: out_word = 8'hED;
		16'hEB12: out_word = 8'hCD;
		16'hEB13: out_word = 8'h95;
		16'hEB14: out_word = 8'h25;
		16'hEB15: out_word = 8'h8F;
		16'hEB16: out_word = 8'h64;
		16'hEB17: out_word = 8'hE5;
		16'hEB18: out_word = 8'hD1;
		16'hEB19: out_word = 8'h5F;
		16'hEB1A: out_word = 8'hB6;
		16'hEB1B: out_word = 8'hE6;
		16'hEB1C: out_word = 8'h7A;
		16'hEB1D: out_word = 8'hB3;
		16'hEB1E: out_word = 8'hB0;
		16'hEB1F: out_word = 8'h7A;
		16'hEB20: out_word = 8'h0F;
		16'hEB21: out_word = 8'hDB;
		16'hEB22: out_word = 8'hFA;
		16'hEB23: out_word = 8'hA1;
		16'hEB24: out_word = 8'h38;
		16'hEB25: out_word = 8'h05;
		16'hEB26: out_word = 8'h7B;
		16'hEB27: out_word = 8'hED;
		16'hEB28: out_word = 8'h18;
		16'hEB29: out_word = 8'hF1;
		16'hEB2A: out_word = 8'h01;
		16'hEB2B: out_word = 8'hFF;
		16'hEB2C: out_word = 8'hBE;
		16'hEB2D: out_word = 8'h9B;
		16'hEB2E: out_word = 8'h2C;
		16'hEB2F: out_word = 8'h3E;
		16'hEB30: out_word = 8'h5F;
		16'hEB31: out_word = 8'hF1;
		16'hEB32: out_word = 8'hC9;
		16'hEB33: out_word = 8'h7E;
		16'hEB34: out_word = 8'hFE;
		16'hEB35: out_word = 8'hE1;
		16'hEB36: out_word = 8'h2E;
		16'hEB37: out_word = 8'hC0;
		16'hEB38: out_word = 8'h23;
		16'hEB39: out_word = 8'hC2;
		16'hEB3A: out_word = 8'h2B;
		16'hEB3B: out_word = 8'h85;
		16'hEB3C: out_word = 8'h20;
		16'hEB3D: out_word = 8'hAF;
		16'hEB3E: out_word = 8'h6E;
		16'hEB3F: out_word = 8'hF4;
		16'hEB40: out_word = 8'h09;
		16'hEB41: out_word = 8'h03;
		16'hEB42: out_word = 8'hF4;
		16'hEB43: out_word = 8'hFD;
		16'hEB44: out_word = 8'h08;
		16'hEB45: out_word = 8'hD0;
		16'hEB46: out_word = 8'h87;
		16'hEB47: out_word = 8'h11;
		16'hEB48: out_word = 8'h8C;
		16'hEB49: out_word = 8'h93;
		16'hEB4A: out_word = 8'h1F;
		16'hEB4B: out_word = 8'hA8;
		16'hEB4C: out_word = 8'h8F;
		16'hEB4D: out_word = 8'h50;
		16'hEB4E: out_word = 8'hE9;
		16'hEB4F: out_word = 8'h9C;
		16'hEB50: out_word = 8'h93;
		16'hEB51: out_word = 8'hA3;
		16'hEB52: out_word = 8'h18;
		16'hEB53: out_word = 8'hC2;
		16'hEB54: out_word = 8'hD0;
		16'hEB55: out_word = 8'hAA;
		16'hEB56: out_word = 8'h81;
		16'hEB57: out_word = 8'hB5;
		16'hEB58: out_word = 8'hC0;
		16'hEB59: out_word = 8'h02;
		16'hEB5A: out_word = 8'h17;
		16'hEB5B: out_word = 8'h04;
		16'hEB5C: out_word = 8'h1C;
		16'hEB5D: out_word = 8'h69;
		16'hEB5E: out_word = 8'h2A;
		16'hEB5F: out_word = 8'h21;
		16'hEB60: out_word = 8'hC5;
		16'hEB61: out_word = 8'h22;
		16'hEB62: out_word = 8'h3B;
		16'hEB63: out_word = 8'h82;
		16'hEB64: out_word = 8'hC9;
		16'hEB65: out_word = 8'h21;
		16'hEB66: out_word = 8'hF9;
		16'hEB67: out_word = 8'h20;
		16'hEB68: out_word = 8'hF6;
		16'hEB69: out_word = 8'hFF;
		16'hEB6A: out_word = 8'h78;
		16'hEB6B: out_word = 8'hA7;
		16'hEB6C: out_word = 8'hC8;
		16'hEB6D: out_word = 8'hC5;
		16'hEB6E: out_word = 8'hCD;
		16'hEB6F: out_word = 8'h71;
		16'hEB70: out_word = 8'h94;
		16'hEB71: out_word = 8'hED;
		16'hEB72: out_word = 8'hC1;
		16'hEB73: out_word = 8'h10;
		16'hEB74: out_word = 8'hF9;
		16'hEB75: out_word = 8'h17;
		16'hEB76: out_word = 8'hF5;
		16'hEB77: out_word = 8'h52;
		16'hEB78: out_word = 8'h93;
		16'hEB79: out_word = 8'hF5;
		16'hEB7A: out_word = 8'h3E;
		16'hEB7B: out_word = 8'hC5;
		16'hEB7C: out_word = 8'hD9;
		16'hEB7D: out_word = 8'h8C;
		16'hEB7E: out_word = 8'hC1;
		16'hEB7F: out_word = 8'h9D;
		16'hEB80: out_word = 8'h05;
		16'hEB81: out_word = 8'h11;
		16'hEB82: out_word = 8'h20;
		16'hEB83: out_word = 8'h00;
		16'hEB84: out_word = 8'h03;
		16'hEB85: out_word = 8'hA3;
		16'hEB86: out_word = 8'hBC;
		16'hEB87: out_word = 8'h0D;
		16'hEB88: out_word = 8'hA2;
		16'hEB89: out_word = 8'h7C;
		16'hEB8A: out_word = 8'h44;
		16'hEB8B: out_word = 8'h03;
		16'hEB8C: out_word = 8'h19;
		16'hEB8D: out_word = 8'h18;
		16'hEB8E: out_word = 8'hF0;
		16'hEB8F: out_word = 8'hF2;
		16'hEB90: out_word = 8'hFC;
		16'hEB91: out_word = 8'h7C;
		16'hEB92: out_word = 8'hFE;
		16'hEB93: out_word = 8'hD2;
		16'hEB94: out_word = 8'hEE;
		16'hEB95: out_word = 8'h95;
		16'hEB96: out_word = 8'hE3;
		16'hEB97: out_word = 8'h16;
		16'hEB98: out_word = 8'h53;
		16'hEB99: out_word = 8'h0F;
		16'hEB9A: out_word = 8'h68;
		16'hEB9B: out_word = 8'h0F;
		16'hEB9C: out_word = 8'h9F;
		16'hEB9D: out_word = 8'h94;
		16'hEB9E: out_word = 8'h32;
		16'hEB9F: out_word = 8'h1E;
		16'hEBA0: out_word = 8'h0B;
		16'hEBA1: out_word = 8'h19;
		16'hEBA2: out_word = 8'h7E;
		16'hEBA3: out_word = 8'hE0;
		16'hEBA4: out_word = 8'hA7;
		16'hEBA5: out_word = 8'hED;
		16'hEBA6: out_word = 8'h52;
		16'hEBA7: out_word = 8'hFC;
		16'hEBA8: out_word = 8'h20;
		16'hEBA9: out_word = 8'hFE;
		16'hEBAA: out_word = 8'h0F;
		16'hEBAB: out_word = 8'h28;
		16'hEBAC: out_word = 8'hDF;
		16'hEBAD: out_word = 8'h89;
		16'hEBAE: out_word = 8'h7E;
		16'hEBAF: out_word = 8'hDB;
		16'hEBB0: out_word = 8'h30;
		16'hEBB1: out_word = 8'hCB;
		16'hEBB2: out_word = 8'hE5;
		16'hEBB3: out_word = 8'hE9;
		16'hEBB4: out_word = 8'hD6;
		16'hEBB5: out_word = 8'hE2;
		16'hEBB6: out_word = 8'hD9;
		16'hEBB7: out_word = 8'h8D;
		16'hEBB8: out_word = 8'h03;
		16'hEBB9: out_word = 8'h18;
		16'hEBBA: out_word = 8'hEB;
		16'hEBBB: out_word = 8'hCE;
		16'hEBBC: out_word = 8'h50;
		16'hEBBD: out_word = 8'h59;
		16'hEBBE: out_word = 8'hC5;
		16'hEBBF: out_word = 8'h82;
		16'hEBC0: out_word = 8'h26;
		16'hEBC1: out_word = 8'h7C;
		16'hEBC2: out_word = 8'h17;
		16'hEBC3: out_word = 8'hBF;
		16'hEBC4: out_word = 8'h8E;
		16'hEBC5: out_word = 8'hE1;
		16'hEBC6: out_word = 8'hA0;
		16'hEBC7: out_word = 8'hA5;
		16'hEBC8: out_word = 8'hC3;
		16'hEBC9: out_word = 8'hF8;
		16'hEBCA: out_word = 8'h7D;
		16'hEBCB: out_word = 8'hAF;
		16'hEBCC: out_word = 8'h23;
		16'hEBCD: out_word = 8'h5B;
		16'hEBCE: out_word = 8'h11;
		16'hEBCF: out_word = 8'h5B;
		16'hEBD0: out_word = 8'hD0;
		16'hEBD1: out_word = 8'hFC;
		16'hEBD2: out_word = 8'hAD;
		16'hEBD3: out_word = 8'h9D;
		16'hEBD4: out_word = 8'hBC;
		16'hEBD5: out_word = 8'hBD;
		16'hEBD6: out_word = 8'h5E;
		16'hEBD7: out_word = 8'hA7;
		16'hEBD8: out_word = 8'hC7;
		16'hEBD9: out_word = 8'h82;
		16'hEBDA: out_word = 8'h10;
		16'hEBDB: out_word = 8'hD6;
		16'hEBDC: out_word = 8'hDC;
		16'hEBDD: out_word = 8'h5F;
		16'hEBDE: out_word = 8'h64;
		16'hEBDF: out_word = 8'h93;
		16'hEBE0: out_word = 8'h28;
		16'hEBE1: out_word = 8'h09;
		16'hEBE2: out_word = 8'h9D;
		16'hEBE3: out_word = 8'h7E;
		16'hEBE4: out_word = 8'h68;
		16'hEBE5: out_word = 8'h18;
		16'hEBE6: out_word = 8'h05;
		16'hEBE7: out_word = 8'hCF;
		16'hEBE8: out_word = 8'hCA;
		16'hEBE9: out_word = 8'h03;
		16'hEBEA: out_word = 8'hCD;
		16'hEBEB: out_word = 8'h21;
		16'hEBEC: out_word = 8'h94;
		16'hEBED: out_word = 8'hE9;
		16'hEBEE: out_word = 8'hFE;
		16'hEBEF: out_word = 8'hFF;
		16'hEBF0: out_word = 8'hC8;
		16'hEBF1: out_word = 8'h9D;
		16'hEBF2: out_word = 8'hF5;
		16'hEBF3: out_word = 8'h4C;
		16'hEBF4: out_word = 8'h9D;
		16'hEBF5: out_word = 8'hF1;
		16'hEBF6: out_word = 8'h7B;
		16'hEBF7: out_word = 8'hA5;
		16'hEBF8: out_word = 8'hE8;
		16'hEBF9: out_word = 8'h9B;
		16'hEBFA: out_word = 8'hEA;
		16'hEBFB: out_word = 8'hB9;
		16'hEBFC: out_word = 8'hAB;
		16'hEBFD: out_word = 8'h17;
		16'hEBFE: out_word = 8'hE2;
		16'hEBFF: out_word = 8'hF4;
		16'hEC00: out_word = 8'h72;
		16'hEC01: out_word = 8'hC8;
		16'hEC02: out_word = 8'h0B;
		16'hEC03: out_word = 8'hF8;
		16'hEC04: out_word = 8'h4A;
		16'hEC05: out_word = 8'hDD;
		16'hEC06: out_word = 8'hF8;
		16'hEC07: out_word = 8'h69;
		16'hEC08: out_word = 8'hDD;
		16'hEC09: out_word = 8'hF4;
		16'hEC0A: out_word = 8'h7B;
		16'hEC0B: out_word = 8'hDF;
		16'hEC0C: out_word = 8'hEF;
		16'hEC0D: out_word = 8'h79;
		16'hEC0E: out_word = 8'hDF;
		16'hEC0F: out_word = 8'hDB;
		16'hEC10: out_word = 8'h3C;
		16'hEC11: out_word = 8'h75;
		16'hEC12: out_word = 8'h2E;
		16'hEC13: out_word = 8'hD5;
		16'hEC14: out_word = 8'hC9;
		16'hEC15: out_word = 8'hF2;
		16'hEC16: out_word = 8'h37;
		16'hEC17: out_word = 8'hF1;
		16'hEC18: out_word = 8'hF9;
		16'hEC19: out_word = 8'hF7;
		16'hEC1A: out_word = 8'h5B;
		16'hEC1B: out_word = 8'hE5;
		16'hEC1C: out_word = 8'hE2;
		16'hEC1D: out_word = 8'h22;
		16'hEC1E: out_word = 8'h31;
		16'hEC1F: out_word = 8'hD7;
		16'hEC20: out_word = 8'hC5;
		16'hEC21: out_word = 8'h33;
		16'hEC22: out_word = 8'h3C;
		16'hEC23: out_word = 8'h3F;
		16'hEC24: out_word = 8'h87;
		16'hEC25: out_word = 8'h02;
		16'hEC26: out_word = 8'h32;
		16'hEC27: out_word = 8'h60;
		16'hEC28: out_word = 8'h6F;
		16'hEC29: out_word = 8'h5A;
		16'hEC2A: out_word = 8'hF9;
		16'hEC2B: out_word = 8'h23;
		16'hEC2C: out_word = 8'h78;
		16'hEC2D: out_word = 8'h96;
		16'hEC2E: out_word = 8'h23;
		16'hEC2F: out_word = 8'hFF;
		16'hEC30: out_word = 8'hAE;
		16'hEC31: out_word = 8'hDC;
		16'hEC32: out_word = 8'hED;
		16'hEC33: out_word = 8'h53;
		16'hEC34: out_word = 8'h11;
		16'hEC35: out_word = 8'hBD;
		16'hEC36: out_word = 8'hE9;
		16'hEC37: out_word = 8'h13;
		16'hEC38: out_word = 8'h11;
		16'hEC39: out_word = 8'h7F;
		16'hEC3A: out_word = 8'h69;
		16'hEC3B: out_word = 8'hE5;
		16'hEC3C: out_word = 8'hDD;
		16'hEC3D: out_word = 8'hAF;
		16'hEC3E: out_word = 8'hE1;
		16'hEC3F: out_word = 8'h87;
		16'hEC40: out_word = 8'h5C;
		16'hEC41: out_word = 8'h5E;
		16'hEC42: out_word = 8'h81;
		16'hEC43: out_word = 8'h16;
		16'hEC44: out_word = 8'h56;
		16'hEC45: out_word = 8'hAB;
		16'hEC46: out_word = 8'h17;
		16'hEC47: out_word = 8'h4C;
		16'hEC48: out_word = 8'h80;
		16'hEC49: out_word = 8'h0C;
		16'hEC4A: out_word = 8'hF6;
		16'hEC4B: out_word = 8'h24;
		16'hEC4C: out_word = 8'hC2;
		16'hEC4D: out_word = 8'hF6;
		16'hEC4E: out_word = 8'h25;
		16'hEC4F: out_word = 8'hC2;
		16'hEC50: out_word = 8'h6E;
		16'hEC51: out_word = 8'h26;
		16'hEC52: out_word = 8'hF5;
		16'hEC53: out_word = 8'h66;
		16'hEC54: out_word = 8'h27;
		16'hEC55: out_word = 8'h22;
		16'hEC56: out_word = 8'h0D;
		16'hEC57: out_word = 8'hE8;
		16'hEC58: out_word = 8'hBF;
		16'hEC59: out_word = 8'h0B;
		16'hEC5A: out_word = 8'h8F;
		16'hEC5B: out_word = 8'h4D;
		16'hEC5C: out_word = 8'hE0;
		16'hEC5D: out_word = 8'h13;
		16'hEC5E: out_word = 8'hEA;
		16'hEC5F: out_word = 8'h14;
		16'hEC60: out_word = 8'hA0;
		16'hEC61: out_word = 8'hE0;
		16'hEC62: out_word = 8'h43;
		16'hEC63: out_word = 8'hF6;
		16'hEC64: out_word = 8'h21;
		16'hEC65: out_word = 8'h33;
		16'hEC66: out_word = 8'hE0;
		16'hEC67: out_word = 8'h22;
		16'hEC68: out_word = 8'hE0;
		16'hEC69: out_word = 8'h23;
		16'hEC6A: out_word = 8'h12;
		16'hEC6B: out_word = 8'h1B;
		16'hEC6C: out_word = 8'h91;
		16'hEC6D: out_word = 8'hE0;
		16'hEC6E: out_word = 8'h19;
		16'hEC6F: out_word = 8'h0C;
		16'hEC70: out_word = 8'hED;
		16'hEC71: out_word = 8'h11;
		16'hEC72: out_word = 8'hCE;
		16'hEC73: out_word = 8'hED;
		16'hEC74: out_word = 8'h12;
		16'hEC75: out_word = 8'hF6;
		16'hEC76: out_word = 8'h09;
		16'hEC77: out_word = 8'hD7;
		16'hEC78: out_word = 8'h9A;
		16'hEC79: out_word = 8'h20;
		16'hEC7A: out_word = 8'h60;
		16'hEC7B: out_word = 8'h69;
		16'hEC7C: out_word = 8'hDD;
		16'hEC7D: out_word = 8'hAA;
		16'hEC7E: out_word = 8'h06;
		16'hEC7F: out_word = 8'hFE;
		16'hEC80: out_word = 8'hDA;
		16'hEC81: out_word = 8'h98;
		16'hEC82: out_word = 8'hEB;
		16'hEC83: out_word = 8'hA4;
		16'hEC84: out_word = 8'h7E;
		16'hEC85: out_word = 8'h19;
		16'hEC86: out_word = 8'h32;
		16'hEC87: out_word = 8'h03;
		16'hEC88: out_word = 8'hDC;
		16'hEC89: out_word = 8'h99;
		16'hEC8A: out_word = 8'h5B;
		16'hEC8B: out_word = 8'hBC;
		16'hEC8C: out_word = 8'h2A;
		16'hEC8D: out_word = 8'hB5;
		16'hEC8E: out_word = 8'hBF;
		16'hEC8F: out_word = 8'h3D;
		16'hEC90: out_word = 8'h21;
		16'hEC91: out_word = 8'h45;
		16'hEC92: out_word = 8'h7F;
		16'hEC93: out_word = 8'h20;
		16'hEC94: out_word = 8'hF8;
		16'hEC95: out_word = 8'hC1;
		16'hEC96: out_word = 8'hCD;
		16'hEC97: out_word = 8'hCE;
		16'hEC98: out_word = 8'h97;
		16'hEC99: out_word = 8'hDD;
		16'hEC9A: out_word = 8'hC5;
		16'hEC9B: out_word = 8'h4E;
		16'hEC9C: out_word = 8'h0E;
		16'hEC9D: out_word = 8'hC8;
		16'hEC9E: out_word = 8'h46;
		16'hEC9F: out_word = 8'h0F;
		16'hECA0: out_word = 8'h7C;
		16'hECA1: out_word = 8'hB4;
		16'hECA2: out_word = 8'hD7;
		16'hECA3: out_word = 8'hF3;
		16'hECA4: out_word = 8'h33;
		16'hECA5: out_word = 8'hC5;
		16'hECA6: out_word = 8'h15;
		16'hECA7: out_word = 8'h51;
		16'hECA8: out_word = 8'h17;
		16'hECA9: out_word = 8'h17;
		16'hECAA: out_word = 8'h44;
		16'hECAB: out_word = 8'h4D;
		16'hECAC: out_word = 8'hCE;
		16'hECAD: out_word = 8'h21;
		16'hECAE: out_word = 8'h19;
		16'hECAF: out_word = 8'hF1;
		16'hECB0: out_word = 8'hAE;
		16'hECB1: out_word = 8'h97;
		16'hECB2: out_word = 8'h7C;
		16'hECB3: out_word = 8'hCA;
		16'hECB4: out_word = 8'h0D;
		16'hECB5: out_word = 8'h32;
		16'hECB6: out_word = 8'h04;
		16'hECB7: out_word = 8'hD7;
		16'hECB8: out_word = 8'hA5;
		16'hECB9: out_word = 8'hBF;
		16'hECBA: out_word = 8'hE8;
		16'hECBB: out_word = 8'h1D;
		16'hECBC: out_word = 8'h22;
		16'hECBD: out_word = 8'h59;
		16'hECBE: out_word = 8'h1F;
		16'hECBF: out_word = 8'h4F;
		16'hECC0: out_word = 8'h3A;
		16'hECC1: out_word = 8'h3C;
		16'hECC2: out_word = 8'hFE;
		16'hECC3: out_word = 8'hFF;
		16'hECC4: out_word = 8'h20;
		16'hECC5: out_word = 8'hE8;
		16'hECC6: out_word = 8'h2B;
		16'hECC7: out_word = 8'h2A;
		16'hECC8: out_word = 8'h1D;
		16'hECC9: out_word = 8'hB5;
		16'hECCA: out_word = 8'h77;
		16'hECCB: out_word = 8'hF2;
		16'hECCC: out_word = 8'hE5;
		16'hECCD: out_word = 8'hD5;
		16'hECCE: out_word = 8'h17;
		16'hECCF: out_word = 8'hB8;
		16'hECD0: out_word = 8'hBF;
		16'hECD1: out_word = 8'hAC;
		16'hECD2: out_word = 8'hF3;
		16'hECD3: out_word = 8'h95;
		16'hECD4: out_word = 8'h3E;
		16'hECD5: out_word = 8'h01;
		16'hECD6: out_word = 8'hD1;
		16'hECD7: out_word = 8'hE1;
		16'hECD8: out_word = 8'hDC;
		16'hECD9: out_word = 8'h28;
		16'hECDA: out_word = 8'h13;
		16'hECDB: out_word = 8'hF1;
		16'hECDC: out_word = 8'h15;
		16'hECDD: out_word = 8'h90;
		16'hECDE: out_word = 8'hEC;
		16'hECDF: out_word = 8'hF4;
		16'hECE0: out_word = 8'h02;
		16'hECE1: out_word = 8'h28;
		16'hECE2: out_word = 8'h01;
		16'hECE3: out_word = 8'hAF;
		16'hECE4: out_word = 8'h0A;
		16'hECE5: out_word = 8'hDF;
		16'hECE6: out_word = 8'hF5;
		16'hECE7: out_word = 8'hA7;
		16'hECE8: out_word = 8'h35;
		16'hECE9: out_word = 8'h0B;
		16'hECEA: out_word = 8'h41;
		16'hECEB: out_word = 8'h5B;
		16'hECEC: out_word = 8'h52;
		16'hECED: out_word = 8'h4B;
		16'hECEE: out_word = 8'h2C;
		16'hECEF: out_word = 8'h66;
		16'hECF0: out_word = 8'h5E;
		16'hECF1: out_word = 8'h2D;
		16'hECF2: out_word = 8'h8C;
		16'hECF3: out_word = 8'h2E;
		16'hECF4: out_word = 8'h66;
		16'hECF5: out_word = 8'h8C;
		16'hECF6: out_word = 8'h2F;
		16'hECF7: out_word = 8'hAB;
		16'hECF8: out_word = 8'h05;
		16'hECF9: out_word = 8'h8C;
		16'hECFA: out_word = 8'hAB;
		16'hECFB: out_word = 8'h8E;
		16'hECFC: out_word = 8'hE6;
		16'hECFD: out_word = 8'hE5;
		16'hECFE: out_word = 8'hD5;
		16'hECFF: out_word = 8'hC5;
		16'hED00: out_word = 8'hAB;
		16'hED01: out_word = 8'h0F;
		16'hED02: out_word = 8'hE6;
		16'hED03: out_word = 8'h46;
		16'hED04: out_word = 8'h21;
		16'hED05: out_word = 8'h11;
		16'hED06: out_word = 8'h68;
		16'hED07: out_word = 8'h8C;
		16'hED08: out_word = 8'hBE;
		16'hED09: out_word = 8'h8C;
		16'hED0A: out_word = 8'h02;
		16'hED0B: out_word = 8'h44;
		16'hED0C: out_word = 8'hE9;
		16'hED0D: out_word = 8'h23;
		16'hED0E: out_word = 8'h30;
		16'hED0F: out_word = 8'hBD;
		16'hED10: out_word = 8'h3E;
		16'hED11: out_word = 8'h3F;
		16'hED12: out_word = 8'hC1;
		16'hED13: out_word = 8'hD1;
		16'hED14: out_word = 8'hF1;
		16'hED15: out_word = 8'hC3;
		16'hED16: out_word = 8'h3D;
		16'hED17: out_word = 8'h93;
		16'hED18: out_word = 8'hFB;
		16'hED19: out_word = 8'hCD;
		16'hED1A: out_word = 8'h99;
		16'hED1B: out_word = 8'h97;
		16'hED1C: out_word = 8'h21;
		16'hED1D: out_word = 8'h0B;
		16'hED1E: out_word = 8'h9F;
		16'hED1F: out_word = 8'h68;
		16'hED20: out_word = 8'h7B;
		16'hED21: out_word = 8'hE6;
		16'hED22: out_word = 8'hF0;
		16'hED23: out_word = 8'hB2;
		16'hED24: out_word = 8'hB1;
		16'hED25: out_word = 8'hEF;
		16'hED26: out_word = 8'hB0;
		16'hED27: out_word = 8'hC9;
		16'hED28: out_word = 8'hD1;
		16'hED29: out_word = 8'h87;
		16'hED2A: out_word = 8'h21;
		16'hED2B: out_word = 8'h7E;
		16'hED2C: out_word = 8'hFE;
		16'hED2D: out_word = 8'h20;
		16'hED2E: out_word = 8'hFC;
		16'hED2F: out_word = 8'h28;
		16'hED30: out_word = 8'h0B;
		16'hED31: out_word = 8'hEB;
		16'hED32: out_word = 8'h36;
		16'hED33: out_word = 8'h2E;
		16'hED34: out_word = 8'h23;
		16'hED35: out_word = 8'h46;
		16'hED36: out_word = 8'h93;
		16'hED37: out_word = 8'hBE;
		16'hED38: out_word = 8'h3E;
		16'hED39: out_word = 8'hF5;
		16'hED3A: out_word = 8'h00;
		16'hED3B: out_word = 8'hE1;
		16'hED3C: out_word = 8'hC9;
		16'hED3D: out_word = 8'hE5;
		16'hED3E: out_word = 8'h3B;
		16'hED3F: out_word = 8'hBB;
		16'hED40: out_word = 8'h36;
		16'hED41: out_word = 8'h43;
		16'hED42: out_word = 8'hF8;
		16'hED43: out_word = 8'h28;
		16'hED44: out_word = 8'hDC;
		16'hED45: out_word = 8'hD9;
		16'hED46: out_word = 8'h0E;
		16'hED47: out_word = 8'h00;
		16'hED48: out_word = 8'hAE;
		16'hED49: out_word = 8'hEE;
		16'hED4A: out_word = 8'h9A;
		16'hED4B: out_word = 8'h7E;
		16'hED4C: out_word = 8'h23;
		16'hED4D: out_word = 8'h08;
		16'hED4E: out_word = 8'h7F;
		16'hED4F: out_word = 8'h71;
		16'hED50: out_word = 8'hE1;
		16'hED51: out_word = 8'h20;
		16'hED52: out_word = 8'h25;
		16'hED53: out_word = 8'h4F;
		16'hED54: out_word = 8'h07;
		16'hED55: out_word = 8'h3E;
		16'hED56: out_word = 8'h05;
		16'hED57: out_word = 8'hFD;
		16'hED58: out_word = 8'hCD;
		16'hED59: out_word = 8'h61;
		16'hED5A: out_word = 8'h96;
		16'hED5B: out_word = 8'hA7;
		16'hED5C: out_word = 8'h28;
		16'hED5D: out_word = 8'h1A;
		16'hED5E: out_word = 8'h7F;
		16'hED5F: out_word = 8'h7B;
		16'hED60: out_word = 8'h3E;
		16'hED61: out_word = 8'h06;
		16'hED62: out_word = 8'h7A;
		16'hED63: out_word = 8'hF5;
		16'hED64: out_word = 8'h0F;
		16'hED65: out_word = 8'h94;
		16'hED66: out_word = 8'hF6;
		16'hED67: out_word = 8'h02;
		16'hED68: out_word = 8'hF6;
		16'hED69: out_word = 8'h77;
		16'hED6A: out_word = 8'hA3;
		16'hED6B: out_word = 8'hB4;
		16'hED6C: out_word = 8'hE5;
		16'hED6D: out_word = 8'h61;
		16'hED6E: out_word = 8'h18;
		16'hED6F: out_word = 8'hD0;
		16'hED70: out_word = 8'h90;
		16'hED71: out_word = 8'hBE;
		16'hED72: out_word = 8'h08;
		16'hED73: out_word = 8'hBD;
		16'hED74: out_word = 8'h50;
		16'hED75: out_word = 8'h47;
		16'hED76: out_word = 8'h2B;
		16'hED77: out_word = 8'h56;
		16'hED78: out_word = 8'hFF;
		16'hED79: out_word = 8'h59;
		16'hED7A: out_word = 8'h7A;
		16'hED7B: out_word = 8'hB3;
		16'hED7C: out_word = 8'hC8;
		16'hED7D: out_word = 8'h7B;
		16'hED7E: out_word = 8'hA7;
		16'hED7F: out_word = 8'hC1;
		16'hED80: out_word = 8'h20;
		16'hED81: out_word = 8'h09;
		16'hED82: out_word = 8'hFF;
		16'hED83: out_word = 8'hFE;
		16'hED84: out_word = 8'h80;
		16'hED85: out_word = 8'h38;
		16'hED86: out_word = 8'h30;
		16'hED87: out_word = 8'h16;
		16'hED88: out_word = 8'h5F;
		16'hED89: out_word = 8'h18;
		16'hED8A: out_word = 8'h2C;
		16'hED8B: out_word = 8'h03;
		16'hED8C: out_word = 8'h04;
		16'hED8D: out_word = 8'h3E;
		16'hED8E: out_word = 8'h0B;
		16'hED8F: out_word = 8'h20;
		16'hED90: out_word = 8'h26;
		16'hED91: out_word = 8'hE7;
		16'hED92: out_word = 8'h7A;
		16'hED93: out_word = 8'h1E;
		16'hED94: out_word = 8'hEF;
		16'hED95: out_word = 8'hF3;
		16'hED96: out_word = 8'hFE;
		16'hED97: out_word = 8'h01;
		16'hED98: out_word = 8'hC0;
		16'hED99: out_word = 8'h28;
		16'hED9A: out_word = 8'h1C;
		16'hED9B: out_word = 8'h85;
		16'hED9C: out_word = 8'hA0;
		16'hED9D: out_word = 8'h51;
		16'hED9E: out_word = 8'h0B;
		16'hED9F: out_word = 8'h16;
		16'hEDA0: out_word = 8'hD6;
		16'hEDA1: out_word = 8'h81;
		16'hEDA2: out_word = 8'h10;
		16'hEDA3: out_word = 8'h80;
		16'hEDA4: out_word = 8'hFC;
		16'hEDA5: out_word = 8'h30;
		16'hEDA6: out_word = 8'h03;
		16'hEDA7: out_word = 8'h7A;
		16'hEDA8: out_word = 8'h18;
		16'hEDA9: out_word = 8'h0E;
		16'hEDAA: out_word = 8'hFE;
		16'hEDAB: out_word = 8'h2F;
		16'hEDAC: out_word = 8'h38;
		16'hEDAD: out_word = 8'h09;
		16'hEDAE: out_word = 8'h1E;
		16'hEDAF: out_word = 8'hB0;
		16'hEDB0: out_word = 8'h0A;
		16'hEDB1: out_word = 8'h40;
		16'hEDB2: out_word = 8'h12;
		16'hEDB3: out_word = 8'h7C;
		16'hEDB4: out_word = 8'hF3;
		16'hEDB5: out_word = 8'h01;
		16'hEDB6: out_word = 8'h83;
		16'hEDB7: out_word = 8'hD9;
		16'hEDB8: out_word = 8'h77;
		16'hEDB9: out_word = 8'h23;
		16'hEDBA: out_word = 8'hF5;
		16'hEDBB: out_word = 8'hAE;
		16'hEDBC: out_word = 8'hC8;
		16'hEDBD: out_word = 8'h18;
		16'hEDBE: out_word = 8'hB8;
		16'hEDBF: out_word = 8'hF3;
		16'hEDC0: out_word = 8'hC9;
		16'hEDC1: out_word = 8'hBD;
		16'hEDC2: out_word = 8'h06;
		16'hEDC3: out_word = 8'hFE;
		16'hEDC4: out_word = 8'h21;
		16'hEDC5: out_word = 8'hF7;
		16'hEDC6: out_word = 8'h0F;
		16'hEDC7: out_word = 8'hED;
		16'hEDC8: out_word = 8'h52;
		16'hEDC9: out_word = 8'hC9;
		16'hEDCA: out_word = 8'h3D;
		16'hEDCB: out_word = 8'hE5;
		16'hEDCC: out_word = 8'hF7;
		16'hEDCD: out_word = 8'hFF;
		16'hEDCE: out_word = 8'h02;
		16'hEDCF: out_word = 8'hF7;
		16'hEDD0: out_word = 8'h0C;
		16'hEDD1: out_word = 8'hED;
		16'hEDD2: out_word = 8'hF1;
		16'hEDD3: out_word = 8'h42;
		16'hEDD4: out_word = 8'hC0;
		16'hEDD5: out_word = 8'h08;
		16'hEDD6: out_word = 8'hF4;
		16'hEDD7: out_word = 8'hDF;
		16'hEDD8: out_word = 8'h71;
		16'hEDD9: out_word = 8'h83;
		16'hEDDA: out_word = 8'h37;
		16'hEDDB: out_word = 8'h3D;
		16'hEDDC: out_word = 8'h6B;
		16'hEDDD: out_word = 8'h18;
		16'hEDDE: out_word = 8'hEF;
		16'hEDDF: out_word = 8'hC2;
		16'hEDE0: out_word = 8'hE9;
		16'hEDE1: out_word = 8'h57;
		16'hEDE2: out_word = 8'hFE;
		16'hEDE3: out_word = 8'hF5;
		16'hEDE4: out_word = 8'h7B;
		16'hEDE5: out_word = 8'h5A;
		16'hEDE6: out_word = 8'h55;
		16'hEDE7: out_word = 8'h4C;
		16'hEDE8: out_word = 8'h9D;
		16'hEDE9: out_word = 8'h86;
		16'hEDEA: out_word = 8'hF4;
		16'hEDEB: out_word = 8'h96;
		16'hEDEC: out_word = 8'hDE;
		16'hEDED: out_word = 8'hD9;
		16'hEDEE: out_word = 8'h77;
		16'hEDEF: out_word = 8'h8F;
		16'hEDF0: out_word = 8'h50;
		16'hEDF1: out_word = 8'hEF;
		16'hEDF2: out_word = 8'h51;
		16'hEDF3: out_word = 8'hF5;
		16'hEDF4: out_word = 8'hC5;
		16'hEDF5: out_word = 8'h8E;
		16'hEDF6: out_word = 8'h21;
		16'hEDF7: out_word = 8'hEF;
		16'hEDF8: out_word = 8'hBB;
		16'hEDF9: out_word = 8'hE5;
		16'hEDFA: out_word = 8'hB5;
		16'hEDFB: out_word = 8'h3B;
		16'hEDFC: out_word = 8'hF1;
		16'hEDFD: out_word = 8'hCB;
		16'hEDFE: out_word = 8'hD6;
		16'hEDFF: out_word = 8'h19;
		16'hEE00: out_word = 8'hBB;
		16'hEE01: out_word = 8'h81;
		16'hEE02: out_word = 8'hC9;
		16'hEE03: out_word = 8'hE0;
		16'hEE04: out_word = 8'h62;
		16'hEE05: out_word = 8'h6B;
		16'hEE06: out_word = 8'h29;
		16'hEE07: out_word = 8'h63;
		16'hEE08: out_word = 8'hCB;
		16'hEE09: out_word = 8'h3C;
		16'hEE0A: out_word = 8'h73;
		16'hEE0B: out_word = 8'h1D;
		16'hEE0C: out_word = 8'h7B;
		16'hEE0D: out_word = 8'h5C;
		16'hEE0E: out_word = 8'hEE;
		16'hEE0F: out_word = 8'h42;
		16'hEE10: out_word = 8'h81;
		16'hEE11: out_word = 8'h4A;
		16'hEE12: out_word = 8'h3B;
		16'hEE13: out_word = 8'hDB;
		16'hEE14: out_word = 8'hF5;
		16'hEE15: out_word = 8'hE5;
		16'hEE16: out_word = 8'h96;
		16'hEE17: out_word = 8'hDA;
		16'hEE18: out_word = 8'h7E;
		16'hEE19: out_word = 8'hE6;
		16'hEE1A: out_word = 8'h01;
		16'hEE1B: out_word = 8'h47;
		16'hEE1C: out_word = 8'h09;
		16'hEE1D: out_word = 8'h46;
		16'hEE1E: out_word = 8'h23;
		16'hEE1F: out_word = 8'hEE;
		16'hEE20: out_word = 8'h83;
		16'hEE21: out_word = 8'hB2;
		16'hEE22: out_word = 8'hC5;
		16'hEE23: out_word = 8'h4B;
		16'hEE24: out_word = 8'hBB;
		16'hEE25: out_word = 8'h13;
		16'hEE26: out_word = 8'hDA;
		16'hEE27: out_word = 8'hC5;
		16'hEE28: out_word = 8'h56;
		16'hEE29: out_word = 8'h58;
		16'hEE2A: out_word = 8'h7C;
		16'hEE2B: out_word = 8'hF5;
		16'hEE2C: out_word = 8'h1F;
		16'hEE2D: out_word = 8'h30;
		16'hEE2E: out_word = 8'h10;
		16'hEE2F: out_word = 8'hCB;
		16'hEE30: out_word = 8'h3A;
		16'hEE31: out_word = 8'h6B;
		16'hEE32: out_word = 8'h1B;
		16'hEE33: out_word = 8'h29;
		16'hEE34: out_word = 8'hFC;
		16'hEE35: out_word = 8'h7A;
		16'hEE36: out_word = 8'hF7;
		16'hEE37: out_word = 8'hE6;
		16'hEE38: out_word = 8'h0F;
		16'hEE39: out_word = 8'h57;
		16'hEE3A: out_word = 8'hC9;
		16'hEE3B: out_word = 8'hF3;
		16'hEE3C: out_word = 8'h48;
		16'hEE3D: out_word = 8'h13;
		16'hEE3E: out_word = 8'hED;
		16'hEE3F: out_word = 8'hD7;
		16'hEE40: out_word = 8'h5B;
		16'hEE41: out_word = 8'h21;
		16'hEE42: out_word = 8'h22;
		16'hEE43: out_word = 8'h48;
		16'hEE44: out_word = 8'h23;
		16'hEE45: out_word = 8'h2F;
		16'hEE46: out_word = 8'hD3;
		16'hEE47: out_word = 8'h8F;
		16'hEE48: out_word = 8'hE5;
		16'hEE49: out_word = 8'hB4;
		16'hEE4A: out_word = 8'hE1;
		16'hEE4B: out_word = 8'hC3;
		16'hEE4C: out_word = 8'h3F;
		16'hEE4D: out_word = 8'hFC;
		16'hEE4E: out_word = 8'h21;
		16'hEE4F: out_word = 8'hFE;
		16'hEE50: out_word = 8'hFF;
		16'hEE51: out_word = 8'hEB;
		16'hEE52: out_word = 8'h19;
		16'hEE53: out_word = 8'h1A;
		16'hEE54: out_word = 8'h23;
		16'hEE55: out_word = 8'h57;
		16'hEE56: out_word = 8'h65;
		16'hEE57: out_word = 8'h3C;
		16'hEE58: out_word = 8'h8D;
		16'hEE59: out_word = 8'h18;
		16'hEE5A: out_word = 8'h08;
		16'hEE5B: out_word = 8'hCB;
		16'hEE5C: out_word = 8'h23;
		16'hEE5D: out_word = 8'h68;
		16'hEE5E: out_word = 8'h12;
		16'hEE5F: out_word = 8'h90;
		16'hEE60: out_word = 8'h15;
		16'hEE61: out_word = 8'hBD;
		16'hEE62: out_word = 8'h14;
		16'hEE63: out_word = 8'h0F;
		16'hEE64: out_word = 8'h30;
		16'hEE65: out_word = 8'hF5;
		16'hEE66: out_word = 8'h79;
		16'hEE67: out_word = 8'hD1;
		16'hEE68: out_word = 8'hFF;
		16'hEE69: out_word = 8'h4E;
		16'hEE6A: out_word = 8'h0A;
		16'hEE6B: out_word = 8'h15;
		16'hEE6C: out_word = 8'h12;
		16'hEE6D: out_word = 8'h1A;
		16'hEE6E: out_word = 8'hD9;
		16'hEE6F: out_word = 8'h59;
		16'hEE70: out_word = 8'h48;
		16'hEE71: out_word = 8'h95;
		16'hEE72: out_word = 8'h04;
		16'hEE73: out_word = 8'h02;
		16'hEE74: out_word = 8'h23;
		16'hEE75: out_word = 8'hDE;
		16'hEE76: out_word = 8'h38;
		16'hEE77: out_word = 8'h19;
		16'hEE78: out_word = 8'h68;
		16'hEE79: out_word = 8'h1A;
		16'hEE7A: out_word = 8'hAA;
		16'hEE7B: out_word = 8'h4F;
		16'hEE7C: out_word = 8'hDE;
		16'hEE7D: out_word = 8'hC9;
		16'hEE7E: out_word = 8'h7E;
		16'hEE7F: out_word = 8'h23;
		16'hEE80: out_word = 8'h93;
		16'hEE81: out_word = 8'h9C;
		16'hEE82: out_word = 8'h5F;
		16'hEE83: out_word = 8'hFC;
		16'hEE84: out_word = 8'h9A;
		16'hEE85: out_word = 8'h57;
		16'hEE86: out_word = 8'hE0;
		16'hEE87: out_word = 8'hFC;
		16'hEE88: out_word = 8'h99;
		16'hEE89: out_word = 8'h4F;
		16'hEE8A: out_word = 8'h69;
		16'hEE8B: out_word = 8'h98;
		16'hEE8C: out_word = 8'h47;
		16'hEE8D: out_word = 8'hF0;
		16'hEE8E: out_word = 8'h83;
		16'hEE8F: out_word = 8'h4A;
		16'hEE90: out_word = 8'hF0;
		16'hEE91: out_word = 8'h8A;
		16'hEE92: out_word = 8'h4C;
		16'hEE93: out_word = 8'hF0;
		16'hEE94: out_word = 8'h89;
		16'hEE95: out_word = 8'hF0;
		16'hEE96: out_word = 8'h88;
		16'hEE97: out_word = 8'hE3;
		16'hEE98: out_word = 8'hF0;
		16'hEE99: out_word = 8'hEB;
		16'hEE9A: out_word = 8'h09;
		16'hEE9B: out_word = 8'h5C;
		16'hEE9C: out_word = 8'h01;
		16'hEE9D: out_word = 8'h08;
		16'hEE9E: out_word = 8'hF0;
		16'hEE9F: out_word = 8'hC9;
		16'hEEA0: out_word = 8'h24;
		16'hEEA1: out_word = 8'h43;
		16'hEEA2: out_word = 8'h20;
		16'hEEA3: out_word = 8'h3C;
		16'hEEA4: out_word = 8'hC5;
		16'hEEA5: out_word = 8'hD5;
		16'hEEA6: out_word = 8'hE5;
		16'hEEA7: out_word = 8'h0E;
		16'hEEA8: out_word = 8'h33;
		16'hEEA9: out_word = 8'hAE;
		16'hEEAA: out_word = 8'h97;
		16'hEEAB: out_word = 8'hFC;
		16'hEEAC: out_word = 8'h1A;
		16'hEEAD: out_word = 8'hA7;
		16'hEEAE: out_word = 8'h28;
		16'hEEAF: out_word = 8'h10;
		16'hEEB0: out_word = 8'h0C;
		16'hEEB1: out_word = 8'hD5;
		16'hEEB2: out_word = 8'hCF;
		16'hEEB3: out_word = 8'h81;
		16'hEEB4: out_word = 8'hFB;
		16'hEEB5: out_word = 8'h81;
		16'hEEB6: out_word = 8'hD1;
		16'hEEB7: out_word = 8'h28;
		16'hEEB8: out_word = 8'h05;
		16'hEEB9: out_word = 8'h51;
		16'hEEBA: out_word = 8'hDA;
		16'hEEBB: out_word = 8'hE6;
		16'hEEBC: out_word = 8'h18;
		16'hEEBD: out_word = 8'hED;
		16'hEEBE: out_word = 8'h79;
		16'hEEBF: out_word = 8'hF6;
		16'hEEC0: out_word = 8'hC1;
		16'hEEC1: out_word = 8'hAD;
		16'hEEC2: out_word = 8'hAA;
		16'hEEC3: out_word = 8'h08;
		16'hEEC4: out_word = 8'h20;
		16'hEEC5: out_word = 8'h05;
		16'hEEC6: out_word = 8'h7F;
		16'hEEC7: out_word = 8'h06;
		16'hEEC8: out_word = 8'h03;
		16'hEEC9: out_word = 8'h1A;
		16'hEECA: out_word = 8'hBE;
		16'hEECB: out_word = 8'hC0;
		16'hEECC: out_word = 8'h23;
		16'hEECD: out_word = 8'h13;
		16'hEECE: out_word = 8'h5C;
		16'hEECF: out_word = 8'hB5;
		16'hEED0: out_word = 8'h5F;
		16'hEED1: out_word = 8'hCE;
		16'hEED2: out_word = 8'hF5;
		16'hEED3: out_word = 8'h22;
		16'hEED4: out_word = 8'h47;
		16'hEED5: out_word = 8'hD7;
		16'hEED6: out_word = 8'hD5;
		16'hEED7: out_word = 8'hF5;
		16'hEED8: out_word = 8'h0E;
		16'hEED9: out_word = 8'hD5;
		16'hEEDA: out_word = 8'h1F;
		16'hEEDB: out_word = 8'hB1;
		16'hEEDC: out_word = 8'hCD;
		16'hEEDD: out_word = 8'h7E;
		16'hEEDE: out_word = 8'hCB;
		16'hEEDF: out_word = 8'h63;
		16'hEEE0: out_word = 8'h28;
		16'hEEE1: out_word = 8'h07;
		16'hEEE2: out_word = 8'hE1;
		16'hEEE3: out_word = 8'hEE;
		16'hEEE4: out_word = 8'hFF;
		16'hEEE5: out_word = 8'h75;
		16'hEEE6: out_word = 8'h18;
		16'hEEE7: out_word = 8'h2A;
		16'hEEE8: out_word = 8'hCD;
		16'hEEE9: out_word = 8'hDB;
		16'hEEEA: out_word = 8'h97;
		16'hEEEB: out_word = 8'hA7;
		16'hEEEC: out_word = 8'hD1;
		16'hEEED: out_word = 8'hEC;
		16'hEEEE: out_word = 8'hCA;
		16'hEEEF: out_word = 8'h5E;
		16'hEEF0: out_word = 8'h98;
		16'hEEF1: out_word = 8'hCD;
		16'hEEF2: out_word = 8'hAD;
		16'hEEF3: out_word = 8'h64;
		16'hEEF4: out_word = 8'hAF;
		16'hEEF5: out_word = 8'hE6;
		16'hEEF6: out_word = 8'hC1;
		16'hEEF7: out_word = 8'hF7;
		16'hEEF8: out_word = 8'hD1;
		16'hEEF9: out_word = 8'hF5;
		16'hEEFA: out_word = 8'h77;
		16'hEEFB: out_word = 8'h98;
		16'hEEFC: out_word = 8'h38;
		16'hEEFD: out_word = 8'h15;
		16'hEEFE: out_word = 8'hCB;
		16'hEEFF: out_word = 8'h53;
		16'hEF00: out_word = 8'hEB;
		16'hEF01: out_word = 8'hBA;
		16'hEF02: out_word = 8'h45;
		16'hEF03: out_word = 8'h1C;
		16'hEF04: out_word = 8'h2A;
		16'hEF05: out_word = 8'h82;
		16'hEF06: out_word = 8'hBC;
		16'hEF07: out_word = 8'h9F;
		16'hEF08: out_word = 8'hB8;
		16'hEF09: out_word = 8'h7A;
		16'hEF0A: out_word = 8'hFE;
		16'hEF0B: out_word = 8'hD0;
		16'hEF0C: out_word = 8'h30;
		16'hEF0D: out_word = 8'h14;
		16'hEF0E: out_word = 8'hA5;
		16'hEF0F: out_word = 8'hD5;
		16'hEF10: out_word = 8'hEA;
		16'hEF11: out_word = 8'hE5;
		16'hEF12: out_word = 8'h71;
		16'hEF13: out_word = 8'h56;
		16'hEF14: out_word = 8'hDD;
		16'hEF15: out_word = 8'h0B;
		16'hEF16: out_word = 8'hC2;
		16'hEF17: out_word = 8'hE1;
		16'hEF18: out_word = 8'hA7;
		16'hEF19: out_word = 8'hF9;
		16'hEF1A: out_word = 8'h42;
		16'hEF1B: out_word = 8'hD1;
		16'hEF1C: out_word = 8'hC2;
		16'hEF1D: out_word = 8'h11;
		16'hEF1E: out_word = 8'h98;
		16'hEF1F: out_word = 8'hF4;
		16'hEF20: out_word = 8'h3F;
		16'hEF21: out_word = 8'hE3;
		16'hEF22: out_word = 8'hC9;
		16'hEF23: out_word = 8'h3A;
		16'hEF24: out_word = 8'h08;
		16'hEF25: out_word = 8'hD0;
		16'hEF26: out_word = 8'hFE;
		16'hEF27: out_word = 8'hF5;
		16'hEF28: out_word = 8'h43;
		16'hEF29: out_word = 8'h37;
		16'hEF2A: out_word = 8'hC0;
		16'hEF2B: out_word = 8'hD5;
		16'hEF2C: out_word = 8'hEF;
		16'hEF2D: out_word = 8'h1E;
		16'hEF2E: out_word = 8'hA7;
		16'hEF2F: out_word = 8'h98;
		16'hEF30: out_word = 8'h0A;
		16'hEF31: out_word = 8'h03;
		16'hEF32: out_word = 8'h8B;
		16'hEF33: out_word = 8'h5F;
		16'hEF34: out_word = 8'h57;
		16'hEF35: out_word = 8'h5C;
		16'hEF36: out_word = 8'h6C;
		16'hEF37: out_word = 8'h9F;
		16'hEF38: out_word = 8'hD1;
		16'hEF39: out_word = 8'hEF;
		16'hEF3A: out_word = 8'hD9;
		16'hEF3B: out_word = 8'h2A;
		16'hEF3C: out_word = 8'h09;
		16'hEF3D: out_word = 8'hD0;
		16'hEF3E: out_word = 8'hAE;
		16'hEF3F: out_word = 8'h2B;
		16'hEF40: out_word = 8'h87;
		16'hEF41: out_word = 8'hA0;
		16'hEF42: out_word = 8'h19;
		16'hEF43: out_word = 8'hDC;
		16'hEF44: out_word = 8'hD9;
		16'hEF45: out_word = 8'hD8;
		16'hEF46: out_word = 8'hF4;
		16'hEF47: out_word = 8'hE9;
		16'hEF48: out_word = 8'h11;
		16'hEF49: out_word = 8'h00;
		16'hEF4A: out_word = 8'h60;
		16'hEF4B: out_word = 8'hE7;
		16'hEF4C: out_word = 8'hD9;
		16'hEF4D: out_word = 8'hE8;
		16'hEF4E: out_word = 8'hC9;
		16'hEF4F: out_word = 8'h3E;
		16'hEF50: out_word = 8'h0F;
		16'hEF51: out_word = 8'h62;
		16'hEF52: out_word = 8'hEC;
		16'hEF53: out_word = 8'hF9;
		16'hEF54: out_word = 8'h81;
		16'hEF55: out_word = 8'h08;
		16'hEF56: out_word = 8'h0A;
		16'hEF57: out_word = 8'h5F;
		16'hEF58: out_word = 8'h57;
		16'hEF59: out_word = 8'hE4;
		16'hEF5A: out_word = 8'hC5;
		16'hEF5B: out_word = 8'h7B;
		16'hEF5C: out_word = 8'h1C;
		16'hEF5D: out_word = 8'h77;
		16'hEF5E: out_word = 8'hFF;
		16'hEF5F: out_word = 8'h48;
		16'hEF60: out_word = 8'h08;
		16'hEF61: out_word = 8'h03;
		16'hEF62: out_word = 8'h3D;
		16'hEF63: out_word = 8'h20;
		16'hEF64: out_word = 8'hEE;
		16'hEF65: out_word = 8'hC9;
		16'hEF66: out_word = 8'hFE;
		16'hEF67: out_word = 8'hF3;
		16'hEF68: out_word = 8'h21;
		16'hEF69: out_word = 8'hFF;
		16'hEF6A: out_word = 8'hF5;
		16'hEF6B: out_word = 8'h22;
		16'hEF6C: out_word = 8'hC8;
		16'hEF6D: out_word = 8'h99;
		16'hEF6E: out_word = 8'h17;
		16'hEF6F: out_word = 8'h55;
		16'hEF70: out_word = 8'h6C;
		16'hEF71: out_word = 8'hCB;
		16'hEF72: out_word = 8'hAE;
		16'hEF73: out_word = 8'hDE;
		16'hEF74: out_word = 8'h7F;
		16'hEF75: out_word = 8'hDE;
		16'hEF76: out_word = 8'h00;
		16'hEF77: out_word = 8'hDA;
		16'hEF78: out_word = 8'hF0;
		16'hEF79: out_word = 8'h75;
		16'hEF7A: out_word = 8'h43;
		16'hEF7B: out_word = 8'hDD;
		16'hEF7C: out_word = 8'h21;
		16'hEF7D: out_word = 8'hC4;
		16'hEF7E: out_word = 8'h7E;
		16'hEF7F: out_word = 8'h66;
		16'hEF80: out_word = 8'hE3;
		16'hEF81: out_word = 8'h73;
		16'hEF82: out_word = 8'h10;
		16'hEF83: out_word = 8'h1C;
		16'hEF84: out_word = 8'hA8;
		16'hEF85: out_word = 8'h56;
		16'hEF86: out_word = 8'hE3;
		16'hEF87: out_word = 8'h11;
		16'hEF88: out_word = 8'h78;
		16'hEF89: out_word = 8'h6B;
		16'hEF8A: out_word = 8'h21;
		16'hEF8B: out_word = 8'h94;
		16'hEF8C: out_word = 8'h66;
		16'hEF8D: out_word = 8'h3E;
		16'hEF8E: out_word = 8'h59;
		16'hEF8F: out_word = 8'h9A;
		16'hEF90: out_word = 8'h01;
		16'hEF91: out_word = 8'h15;
		16'hEF92: out_word = 8'hBD;
		16'hEF93: out_word = 8'h17;
		16'hEF94: out_word = 8'hEB;
		16'hEF95: out_word = 8'h8F;
		16'hEF96: out_word = 8'hD9;
		16'hEF97: out_word = 8'h36;
		16'hEF98: out_word = 8'hC5;
		16'hEF99: out_word = 8'h0D;
		16'hEF9A: out_word = 8'h23;
		16'hEF9B: out_word = 8'h8A;
		16'hEF9C: out_word = 8'h03;
		16'hEF9D: out_word = 8'h05;
		16'hEF9E: out_word = 8'h7E;
		16'hEF9F: out_word = 8'h7A;
		16'hEFA0: out_word = 8'hEC;
		16'hEFA1: out_word = 8'h81;
		16'hEFA2: out_word = 8'h3F;
		16'hEFA3: out_word = 8'hD6;
		16'hEFA4: out_word = 8'h04;
		16'hEFA5: out_word = 8'h87;
		16'hEFA6: out_word = 8'h4F;
		16'hEFA7: out_word = 8'hFF;
		16'hEFA8: out_word = 8'hD9;
		16'hEFA9: out_word = 8'hEB;
		16'hEFAA: out_word = 8'h21;
		16'hEFAB: out_word = 8'h7B;
		16'hEFAC: out_word = 8'hAC;
		16'hEFAD: out_word = 8'h6B;
		16'hEFAE: out_word = 8'hF3;
		16'hEFAF: out_word = 8'h41;
		16'hEFB0: out_word = 8'h09;
		16'hEFB1: out_word = 8'h01;
		16'hEFB2: out_word = 8'h10;
		16'hEFB3: out_word = 8'hD2;
		16'hEFB4: out_word = 8'h7D;
		16'hEFB5: out_word = 8'h1A;
		16'hEFB6: out_word = 8'h0F;
		16'hEFB7: out_word = 8'h7F;
		16'hEFB8: out_word = 8'hFF;
		16'hEFB9: out_word = 8'hE6;
		16'hEFBA: out_word = 8'h1F;
		16'hEFBB: out_word = 8'hC6;
		16'hEFBC: out_word = 8'h45;
		16'hEFBD: out_word = 8'h12;
		16'hEFBE: out_word = 8'h13;
		16'hEFBF: out_word = 8'h24;
		16'hEFC0: out_word = 8'hD0;
		16'hEFC1: out_word = 8'hD9;
		16'hEFC2: out_word = 8'h69;
		16'hEFC3: out_word = 8'h4F;
		16'hEFC4: out_word = 8'hE0;
		16'hEFC5: out_word = 8'hE7;
		16'hEFC6: out_word = 8'h81;
		16'hEFC7: out_word = 8'h21;
		16'hEFC8: out_word = 8'hDB;
		16'hEFC9: out_word = 8'hE1;
		16'hEFCA: out_word = 8'h09;
		16'hEFCB: out_word = 8'h0E;
		16'hEFCC: out_word = 8'hB9;
		16'hEFCD: out_word = 8'h05;
		16'hEFCE: out_word = 8'hC0;
		16'hEFCF: out_word = 8'h19;
		16'hEFD0: out_word = 8'hD7;
		16'hEFD1: out_word = 8'h10;
		16'hEFD2: out_word = 8'hBD;
		16'hEFD3: out_word = 8'hBE;
		16'hEFD4: out_word = 8'h24;
		16'hEFD5: out_word = 8'h23;
		16'hEFD6: out_word = 8'hDD;
		16'hEFD7: out_word = 8'h46;
		16'hEFD8: out_word = 8'h02;
		16'hEFD9: out_word = 8'h05;
		16'hEFDA: out_word = 8'h3F;
		16'hEFDB: out_word = 8'h48;
		16'hEFDC: out_word = 8'h3E;
		16'hEFDD: out_word = 8'h65;
		16'hEFDE: out_word = 8'hA8;
		16'hEFDF: out_word = 8'h70;
		16'hEFE0: out_word = 8'h7F;
		16'hEFE1: out_word = 8'h33;
		16'hEFE2: out_word = 8'h3C;
		16'hEFE3: out_word = 8'h10;
		16'hEFE4: out_word = 8'hFB;
		16'hEFE5: out_word = 8'h22;
		16'hEFE6: out_word = 8'h84;
		16'hEFE7: out_word = 8'h66;
		16'hEFE8: out_word = 8'h41;
		16'hEFE9: out_word = 8'hCC;
		16'hEFEA: out_word = 8'h36;
		16'hEFEB: out_word = 8'h61;
		16'hEFEC: out_word = 8'hA7;
		16'hEFED: out_word = 8'h99;
		16'hEFEE: out_word = 8'h5F;
		16'hEFEF: out_word = 8'h10;
		16'hEFF0: out_word = 8'hF8;
		16'hEFF1: out_word = 8'h79;
		16'hEFF2: out_word = 8'hD9;
		16'hEFF3: out_word = 8'hF8;
		16'hEFF4: out_word = 8'h3D;
		16'hEFF5: out_word = 8'h28;
		16'hEFF6: out_word = 8'h06;
		16'hEFF7: out_word = 8'hCD;
		16'hEFF8: out_word = 8'hB2;
		16'hEFF9: out_word = 8'h3F;
		16'hEFFA: out_word = 8'hC3;
		16'hEFFB: out_word = 8'h83;
		16'hEFFC: out_word = 8'h60;
		16'hEFFD: out_word = 8'hF3;
		16'hEFFE: out_word = 8'hDD;
		16'hEFFF: out_word = 8'hD2;
		16'hF000: out_word = 8'h7E;
		16'hF001: out_word = 8'h12;
		16'hF002: out_word = 8'h6A;
		16'hF003: out_word = 8'h01;
		16'hF004: out_word = 8'hE8;
		16'hF005: out_word = 8'h1A;
		16'hF006: out_word = 8'h1E;
		16'hF007: out_word = 8'h32;
		16'hF008: out_word = 8'hC0;
		16'hF009: out_word = 8'h70;
		16'hF00A: out_word = 8'hF9;
		16'hF00B: out_word = 8'h09;
		16'hF00C: out_word = 8'h21;
		16'hF00D: out_word = 8'h01;
		16'hF00E: out_word = 8'h17;
		16'hF00F: out_word = 8'hF8;
		16'hF010: out_word = 8'hF4;
		16'hF011: out_word = 8'h20;
		16'hF012: out_word = 8'h16;
		16'hF013: out_word = 8'hC5;
		16'hF014: out_word = 8'h77;
		16'hF015: out_word = 8'h4B;
		16'hF016: out_word = 8'hB7;
		16'hF017: out_word = 8'hEF;
		16'hF018: out_word = 8'h01;
		16'hF019: out_word = 8'hC1;
		16'hF01A: out_word = 8'hEF;
		16'hF01B: out_word = 8'hAE;
		16'hF01C: out_word = 8'hE6;
		16'hF01D: out_word = 8'h10;
		16'hF01E: out_word = 8'h4C;
		16'hF01F: out_word = 8'h1C;
		16'hF020: out_word = 8'h28;
		16'hF021: out_word = 8'h11;
		16'hF022: out_word = 8'hFF;
		16'hF023: out_word = 8'h45;
		16'hF024: out_word = 8'hD8;
		16'hF025: out_word = 8'h68;
		16'hF026: out_word = 8'hC3;
		16'hF027: out_word = 8'h2C;
		16'hF028: out_word = 8'h84;
		16'hF029: out_word = 8'hF3;
		16'hF02A: out_word = 8'hCD;
		16'hF02B: out_word = 8'hF8;
		16'hF02C: out_word = 8'h59;
		16'hF02D: out_word = 8'h63;
		16'hF02E: out_word = 8'hDD;
		16'hF02F: out_word = 8'h6E;
		16'hF030: out_word = 8'h12;
		16'hF031: out_word = 8'hBA;
		16'hF032: out_word = 8'h66;
		16'hF033: out_word = 8'h13;
		16'hF034: out_word = 8'h5D;
		16'hF035: out_word = 8'hCA;
		16'hF036: out_word = 8'h29;
		16'hF037: out_word = 8'hF5;
		16'hF038: out_word = 8'h8C;
		16'hF039: out_word = 8'hD2;
		16'hF03A: out_word = 8'h99;
		16'hF03B: out_word = 8'hD4;
		16'hF03C: out_word = 8'h23;
		16'hF03D: out_word = 8'h8D;
		16'hF03E: out_word = 8'hD0;
		16'hF03F: out_word = 8'h76;
		16'hF040: out_word = 8'h7F;
		16'hF041: out_word = 8'h7A;
		16'hF042: out_word = 8'hCF;
		16'hF043: out_word = 8'h28;
		16'hF044: out_word = 8'h4C;
		16'hF045: out_word = 8'hC5;
		16'hF046: out_word = 8'h74;
		16'hF047: out_word = 8'hF0;
		16'hF048: out_word = 8'h02;
		16'hF049: out_word = 8'hC1;
		16'hF04A: out_word = 8'h7A;
		16'hF04B: out_word = 8'hC6;
		16'hF04C: out_word = 8'h5B;
		16'hF04D: out_word = 8'h04;
		16'hF04E: out_word = 8'hEE;
		16'hF04F: out_word = 8'h22;
		16'hF050: out_word = 8'h23;
		16'hF051: out_word = 8'h7E;
		16'hF052: out_word = 8'hDA;
		16'hF053: out_word = 8'hEE;
		16'hF054: out_word = 8'hF9;
		16'hF055: out_word = 8'hF3;
		16'hF056: out_word = 8'h09;
		16'hF057: out_word = 8'h38;
		16'hF058: out_word = 8'hC6;
		16'hF059: out_word = 8'h72;
		16'hF05A: out_word = 8'h13;
		16'hF05B: out_word = 8'h5B;
		16'hF05C: out_word = 8'h77;
		16'hF05D: out_word = 8'h0F;
		16'hF05E: out_word = 8'h57;
		16'hF05F: out_word = 8'h8D;
		16'hF060: out_word = 8'hDD;
		16'hF061: out_word = 8'h71;
		16'hF062: out_word = 8'h10;
		16'hF063: out_word = 8'h17;
		16'hF064: out_word = 8'h70;
		16'hF065: out_word = 8'h11;
		16'hF066: out_word = 8'hE1;
		16'hF067: out_word = 8'hC3;
		16'hF068: out_word = 8'h3E;
		16'hF069: out_word = 8'h84;
		16'hF06A: out_word = 8'h4E;
		16'hF06B: out_word = 8'h56;
		16'hF06C: out_word = 8'hEA;
		16'hF06D: out_word = 8'h5E;
		16'hF06E: out_word = 8'h12;
		16'hF06F: out_word = 8'h7C;
		16'hF070: out_word = 8'h6C;
		16'hF071: out_word = 8'h0F;
		16'hF072: out_word = 8'h72;
		16'hF073: out_word = 8'h2B;
		16'hF074: out_word = 8'h73;
		16'hF075: out_word = 8'h68;
		16'hF076: out_word = 8'h77;
		16'hF077: out_word = 8'h88;
		16'hF078: out_word = 8'hD5;
		16'hF079: out_word = 8'hD4;
		16'hF07A: out_word = 8'hDE;
		16'hF07B: out_word = 8'h8C;
		16'hF07C: out_word = 8'h8D;
		16'hF07D: out_word = 8'hBF;
		16'hF07E: out_word = 8'hF5;
		16'hF07F: out_word = 8'h24;
		16'hF080: out_word = 8'hED;
		16'hF081: out_word = 8'h53;
		16'hF082: out_word = 8'h49;
		16'hF083: out_word = 8'hCB;
		16'hF084: out_word = 8'hC8;
		16'hF085: out_word = 8'h4B;
		16'hF086: out_word = 8'hF7;
		16'hF087: out_word = 8'h8C;
		16'hF088: out_word = 8'h7A;
		16'hF089: out_word = 8'h5F;
		16'hF08A: out_word = 8'hDF;
		16'hF08B: out_word = 8'h77;
		16'hF08C: out_word = 8'hFC;
		16'hF08D: out_word = 8'hE4;
		16'hF08E: out_word = 8'h7E;
		16'hF08F: out_word = 8'hD6;
		16'hF090: out_word = 8'h04;
		16'hF091: out_word = 8'h08;
		16'hF092: out_word = 8'h8A;
		16'hF093: out_word = 8'h9D;
		16'hF094: out_word = 8'h78;
		16'hF095: out_word = 8'h93;
		16'hF096: out_word = 8'h58;
		16'hF097: out_word = 8'h11;
		16'hF098: out_word = 8'h01;
		16'hF099: out_word = 8'hA3;
		16'hF09A: out_word = 8'h7C;
		16'hF09B: out_word = 8'hFF;
		16'hF09C: out_word = 8'h02;
		16'hF09D: out_word = 8'h75;
		16'hF09E: out_word = 8'hED;
		16'hF09F: out_word = 8'hB0;
		16'hF0A0: out_word = 8'hCF;
		16'hF0A1: out_word = 8'hF4;
		16'hF0A2: out_word = 8'hD7;
		16'hF0A3: out_word = 8'hBF;
		16'hF0A4: out_word = 8'h42;
		16'hF0A5: out_word = 8'h06;
		16'hF0A6: out_word = 8'h01;
		16'hF0A7: out_word = 8'h3E;
		16'hF0A8: out_word = 8'hF6;
		16'hF0A9: out_word = 8'hD5;
		16'hF0AA: out_word = 8'h21;
		16'hF0AB: out_word = 8'hD0;
		16'hF0AC: out_word = 8'h70;
		16'hF0AD: out_word = 8'h0E;
		16'hF0AE: out_word = 8'h5E;
		16'hF0AF: out_word = 8'h04;
		16'hF0B0: out_word = 8'h7F;
		16'hF0B1: out_word = 8'hF7;
		16'hF0B2: out_word = 8'hF5;
		16'hF0B3: out_word = 8'hCD;
		16'hF0B4: out_word = 8'h8F;
		16'hF0B5: out_word = 8'h62;
		16'hF0B6: out_word = 8'hF1;
		16'hF0B7: out_word = 8'hC9;
		16'hF0B8: out_word = 8'h60;
		16'hF0B9: out_word = 8'h10;
		16'hF0BA: out_word = 8'h00;
		16'hF0BB: out_word = 8'hFC;
		16'hF0BC: out_word = 8'h78;
		16'hF0BD: out_word = 8'h84;
		16'hF0BE: out_word = 8'h9F;
		16'hF0BF: out_word = 8'hA1;
		16'hF0C0: out_word = 8'hC2;
		16'hF0C1: out_word = 8'hFC;
		16'hF0C2: out_word = 8'h10;
		16'hF0C3: out_word = 8'h23;
		16'hF0C4: out_word = 8'hFE;
		16'hF0C5: out_word = 8'hC8;
		16'hF0C6: out_word = 8'h82;
		16'hF0C7: out_word = 8'hFF;
		16'hF0C8: out_word = 8'h60;
		16'hF0C9: out_word = 8'h71;
		16'hF0CA: out_word = 8'h38;
		16'hF0CB: out_word = 8'h7C;
		16'hF0CC: out_word = 8'h54;
		16'hF0CD: out_word = 8'hB0;
		16'hF0CE: out_word = 8'h44;
		16'hF0CF: out_word = 8'h6C;
		16'hF0D0: out_word = 8'hC1;
		16'hF0D1: out_word = 8'hC9;
		16'hF0D2: out_word = 8'h00;
		16'hF0D3: out_word = 8'h28;
		16'hF0D4: out_word = 8'hFB;
		16'hF0D5: out_word = 8'hFA;
		16'hF0D6: out_word = 8'h91;
		16'hF0D7: out_word = 8'h10;
		16'hF0D8: out_word = 8'hE8;
		16'hF0D9: out_word = 8'h43;
		16'hF0DA: out_word = 8'h68;
		16'hF0DB: out_word = 8'hF8;
		16'hF0DC: out_word = 8'h24;
		16'hF0DD: out_word = 8'hFC;
		16'hF0DE: out_word = 8'hE7;
		16'hF0DF: out_word = 8'h62;
		16'hF0E0: out_word = 8'hF3;
		16'hF0E1: out_word = 8'hF0;
		16'hF0E2: out_word = 8'hF0;
		16'hF0E3: out_word = 8'hC8;
		16'hF0E4: out_word = 8'hF8;
		16'hF0E5: out_word = 8'h3E;
		16'hF0E6: out_word = 8'h30;
		16'hF0E7: out_word = 8'h78;
		16'hF0E8: out_word = 8'h38;
		16'hF0E9: out_word = 8'hA6;
		16'hF0EA: out_word = 8'hFA;
		16'hF0EB: out_word = 8'hFC;
		16'hF0EC: out_word = 8'h3E;
		16'hF0ED: out_word = 8'hCC;
		16'hF0EE: out_word = 8'h84;
		16'hF0EF: out_word = 8'h38;
		16'hF0F0: out_word = 8'hA5;
		16'hF0F1: out_word = 8'hFA;
		16'hF0F2: out_word = 8'h23;
		16'hF0F3: out_word = 8'hF0;
		16'hF0F4: out_word = 8'h48;
		16'hF0F5: out_word = 8'hB4;
		16'hF0F6: out_word = 8'h47;
		16'hF0F7: out_word = 8'hF0;
		16'hF0F8: out_word = 8'hB4;
		16'hF0F9: out_word = 8'h4E;
		16'hF0FA: out_word = 8'hF0;
		16'hF0FB: out_word = 8'h1C;
		16'hF0FC: out_word = 8'h0C;
		16'hF0FD: out_word = 8'h14;
		16'hF0FE: out_word = 8'hF1;
		16'hF0FF: out_word = 8'hEF;
		16'hF100: out_word = 8'hC8;
		16'hF101: out_word = 8'h8E;
		16'hF102: out_word = 8'h44;
		16'hF103: out_word = 8'h4E;
		16'hF104: out_word = 8'hC5;
		16'hF105: out_word = 8'hFE;
		16'hF106: out_word = 8'h3C;
		16'hF107: out_word = 8'h24;
		16'hF108: out_word = 8'h34;
		16'hF109: out_word = 8'h20;
		16'hF10A: out_word = 8'h7C;
		16'hF10B: out_word = 8'h60;
		16'hF10C: out_word = 8'hE0;
		16'hF10D: out_word = 8'h62;
		16'hF10E: out_word = 8'hA3;
		16'hF10F: out_word = 8'h31;
		16'hF110: out_word = 8'hEF;
		16'hF111: out_word = 8'hE7;
		16'hF112: out_word = 8'h4C;
		16'hF113: out_word = 8'hCC;
		16'hF114: out_word = 8'hC0;
		16'hF115: out_word = 8'hB2;
		16'hF116: out_word = 8'h38;
		16'hF117: out_word = 8'h6C;
		16'hF118: out_word = 8'h1C;
		16'hF119: out_word = 8'h50;
		16'hF11A: out_word = 8'hCF;
		16'hF11B: out_word = 8'hA7;
		16'hF11C: out_word = 8'h40;
		16'hF11D: out_word = 8'h60;
		16'hF11E: out_word = 8'h70;
		16'hF11F: out_word = 8'h8C;
		16'hF120: out_word = 8'h78;
		16'hF121: out_word = 8'h20;
		16'hF122: out_word = 8'h40;
		16'hF123: out_word = 8'h70;
		16'hF124: out_word = 8'h08;
		16'hF125: out_word = 8'h18;
		16'hF126: out_word = 8'h38;
		16'hF127: out_word = 8'h06;
		16'hF128: out_word = 8'h10;
		16'hF129: out_word = 8'h24;
		16'hF12A: out_word = 8'hA1;
		16'hF12B: out_word = 8'h14;
		16'hF12C: out_word = 8'h44;
		16'hF12D: out_word = 8'h8F;
		16'hF12E: out_word = 8'h28;
		16'hF12F: out_word = 8'h80;
		16'hF130: out_word = 8'hFF;
		16'hF131: out_word = 8'h4E;
		16'hF132: out_word = 8'hFB;
		16'hF133: out_word = 8'hC0;
		16'hF134: out_word = 8'h3C;
		16'hF135: out_word = 8'h54;
		16'hF136: out_word = 8'h71;
		16'hF137: out_word = 8'hFF;
		16'hF138: out_word = 8'h34;
		16'hF139: out_word = 8'h14;
		16'hF13A: out_word = 8'hCC;
		16'hF13B: out_word = 8'hB8;
		16'hF13C: out_word = 8'h40;
		16'hF13D: out_word = 8'h8D;
		16'hF13E: out_word = 8'hB0;
		16'hF13F: out_word = 8'h08;
		16'hF140: out_word = 8'h80;
		16'hF141: out_word = 8'h70;
		16'hF142: out_word = 8'hE1;
		16'hF143: out_word = 8'hFF;
		16'hF144: out_word = 8'h86;
		16'hF145: out_word = 8'h71;
		16'hF146: out_word = 8'h79;
		16'hF147: out_word = 8'hC0;
		16'hF148: out_word = 8'hD9;
		16'hF149: out_word = 8'hDE;
		16'hF14A: out_word = 8'hF7;
		16'hF14B: out_word = 8'h05;
		16'hF14C: out_word = 8'hC6;
		16'hF14D: out_word = 8'h58;
		16'hF14E: out_word = 8'h84;
		16'hF14F: out_word = 8'hC9;
		16'hF150: out_word = 8'hF7;
		16'hF151: out_word = 8'h80;
		16'hF152: out_word = 8'h18;
		16'hF153: out_word = 8'h33;
		16'hF154: out_word = 8'hD0;
		16'hF155: out_word = 8'hF8;
		16'hF156: out_word = 8'h30;
		16'hF157: out_word = 8'h06;
		16'hF158: out_word = 8'h70;
		16'hF159: out_word = 8'hF8;
		16'hF15A: out_word = 8'h9A;
		16'hF15B: out_word = 8'h9E;
		16'hF15C: out_word = 8'hFF;
		16'hF15D: out_word = 8'h7C;
		16'hF15E: out_word = 8'h48;
		16'hF15F: out_word = 8'hF9;
		16'hF160: out_word = 8'h48;
		16'hF161: out_word = 8'h6A;
		16'hF162: out_word = 8'hC2;
		16'hF163: out_word = 8'h00;
		16'hF164: out_word = 8'hD0;
		16'hF165: out_word = 8'h2F;
		16'hF166: out_word = 8'hE3;
		16'hF167: out_word = 8'hE9;
		16'hF168: out_word = 8'hCD;
		16'hF169: out_word = 8'h29;
		16'hF16A: out_word = 8'hC8;
		16'hF16B: out_word = 8'hFF;
		16'hF16C: out_word = 8'hC0;
		16'hF16D: out_word = 8'h88;
		16'hF16E: out_word = 8'hBA;
		16'hF16F: out_word = 8'hEF;
		16'hF170: out_word = 8'h8F;
		16'hF171: out_word = 8'h8A;
		16'hF172: out_word = 8'h01;
		16'hF173: out_word = 8'hFF;
		16'hF174: out_word = 8'h7C;
		16'hF175: out_word = 8'h19;
		16'hF176: out_word = 8'h10;
		16'hF177: out_word = 8'hFD;
		16'hF178: out_word = 8'hE8;
		16'hF179: out_word = 8'h08;
		16'hF17A: out_word = 8'h50;
		16'hF17B: out_word = 8'h31;
		16'hF17C: out_word = 8'h14;
		16'hF17D: out_word = 8'h0E;
		16'hF17E: out_word = 8'hE7;
		16'hF17F: out_word = 8'hC4;
		16'hF180: out_word = 8'hC8;
		16'hF181: out_word = 8'h27;
		16'hF182: out_word = 8'h20;
		16'hF183: out_word = 8'h4C;
		16'hF184: out_word = 8'h8C;
		16'hF185: out_word = 8'h48;
		16'hF186: out_word = 8'hF0;
		16'hF187: out_word = 8'h28;
		16'hF188: out_word = 8'h1D;
		16'hF189: out_word = 8'h2C;
		16'hF18A: out_word = 8'h48;
		16'hF18B: out_word = 8'h34;
		16'hF18C: out_word = 8'h2F;
		16'hF18D: out_word = 8'hF8;
		16'hF18E: out_word = 8'h20;
		16'hF18F: out_word = 8'h17;
		16'hF190: out_word = 8'hD9;
		16'hF191: out_word = 8'h48;
		16'hF192: out_word = 8'h03;
		16'hF193: out_word = 8'hC7;
		16'hF194: out_word = 8'h41;
		16'hF195: out_word = 8'hF0;
		16'hF196: out_word = 8'h10;
		16'hF197: out_word = 8'hFF;
		16'hF198: out_word = 8'h37;
		16'hF199: out_word = 8'h09;
		16'hF19A: out_word = 8'hC7;
		16'hF19B: out_word = 8'hCE;
		16'hF19C: out_word = 8'hDC;
		16'hF19D: out_word = 8'h79;
		16'hF19E: out_word = 8'hAF;
		16'hF19F: out_word = 8'h1B;
		16'hF1A0: out_word = 8'h67;
		16'hF1A1: out_word = 8'h2F;
		16'hF1A2: out_word = 8'hA4;
		16'hF1A3: out_word = 8'h20;
		16'hF1A4: out_word = 8'h36;
		16'hF1A5: out_word = 8'h8E;
		16'hF1A6: out_word = 8'h57;
		16'hF1A7: out_word = 8'h94;
		16'hF1A8: out_word = 8'h30;
		16'hF1A9: out_word = 8'hF3;
		16'hF1AA: out_word = 8'hE8;
		16'hF1AB: out_word = 8'h04;
		16'hF1AC: out_word = 8'h08;
		16'hF1AD: out_word = 8'hEB;
		16'hF1AE: out_word = 8'h40;
		16'hF1AF: out_word = 8'hAF;
		16'hF1B0: out_word = 8'h80;
		16'hF1B1: out_word = 8'hCC;
		16'hF1B2: out_word = 8'hE0;
		16'hF1B3: out_word = 8'h4C;
		16'hF1B4: out_word = 8'h20;
		16'hF1B5: out_word = 8'h64;
		16'hF1B6: out_word = 8'h37;
		16'hF1B7: out_word = 8'h10;
		16'hF1B8: out_word = 8'h51;
		16'hF1B9: out_word = 8'hB8;
		16'hF1BA: out_word = 8'h07;
		16'hF1BB: out_word = 8'h7E;
		16'hF1BC: out_word = 8'hD0;
		16'hF1BD: out_word = 8'h04;
		16'hF1BE: out_word = 8'h13;
		16'hF1BF: out_word = 8'h82;
		16'hF1C0: out_word = 8'h50;
		16'hF1C1: out_word = 8'h91;
		16'hF1C2: out_word = 8'hF9;
		16'hF1C3: out_word = 8'hA5;
		16'hF1C4: out_word = 8'h44;
		16'hF1C5: out_word = 8'hF0;
		16'hF1C6: out_word = 8'h7F;
		16'hF1C7: out_word = 8'hE8;
		16'hF1C8: out_word = 8'h28;
		16'hF1C9: out_word = 8'h48;
		16'hF1CA: out_word = 8'h86;
		16'hF1CB: out_word = 8'h7C;
		16'hF1CC: out_word = 8'h9B;
		16'hF1CD: out_word = 8'hF0;
		16'hF1CE: out_word = 8'h40;
		16'hF1CF: out_word = 8'h78;
		16'hF1D0: out_word = 8'hC2;
		16'hF1D1: out_word = 8'hF0;
		16'hF1D2: out_word = 8'h95;
		16'hF1D3: out_word = 8'hF8;
		16'hF1D4: out_word = 8'hF7;
		16'hF1D5: out_word = 8'hAE;
		16'hF1D6: out_word = 8'h1C;
		16'hF1D7: out_word = 8'hE0;
		16'hF1D8: out_word = 8'h86;
		16'hF1D9: out_word = 8'h70;
		16'hF1DA: out_word = 8'hD0;
		16'hF1DB: out_word = 8'h67;
		16'hF1DC: out_word = 8'h92;
		16'hF1DD: out_word = 8'hF0;
		16'hF1DE: out_word = 8'hFA;
		16'hF1DF: out_word = 8'h3C;
		16'hF1E0: out_word = 8'h5E;
		16'hF1E1: out_word = 8'hCD;
		16'hF1E2: out_word = 8'h92;
		16'hF1E3: out_word = 8'h2F;
		16'hF1E4: out_word = 8'hFD;
		16'hF1E5: out_word = 8'h35;
		16'hF1E6: out_word = 8'h00;
		16'hF1E7: out_word = 8'h22;
		16'hF1E8: out_word = 8'h88;
		16'hF1E9: out_word = 8'h98;
		16'hF1EA: out_word = 8'h3C;
		16'hF1EB: out_word = 8'h60;
		16'hF1EC: out_word = 8'h81;
		16'hF1ED: out_word = 8'hF2;
		16'hF1EE: out_word = 8'h7F;
		16'hF1EF: out_word = 8'h22;
		16'hF1F0: out_word = 8'hF2;
		16'hF1F1: out_word = 8'hE9;
		16'hF1F2: out_word = 8'h23;
		16'hF1F3: out_word = 8'hD0;
		16'hF1F4: out_word = 8'h52;
		16'hF1F5: out_word = 8'hD1;
		16'hF1F6: out_word = 8'hC0;
		16'hF1F7: out_word = 8'h5C;
		16'hF1F8: out_word = 8'hEF;
		16'hF1F9: out_word = 8'h40;
		16'hF1FA: out_word = 8'h3B;
		16'hF1FB: out_word = 8'hC0;
		16'hF1FC: out_word = 8'hE4;
		16'hF1FD: out_word = 8'h66;
		16'hF1FE: out_word = 8'hF8;
		16'hF1FF: out_word = 8'hA0;
		16'hF200: out_word = 8'hA2;
		16'hF201: out_word = 8'hA0;
		16'hF202: out_word = 8'h6E;
		16'hF203: out_word = 8'h47;
		16'hF204: out_word = 8'hF0;
		16'hF205: out_word = 8'h40;
		16'hF206: out_word = 8'h71;
		16'hF207: out_word = 8'hA8;
		16'hF208: out_word = 8'h11;
		16'hF209: out_word = 8'hF2;
		16'hF20A: out_word = 8'hF0;
		16'hF20B: out_word = 8'hE5;
		16'hF20C: out_word = 8'h80;
		16'hF20D: out_word = 8'hF6;
		16'hF20E: out_word = 8'hB8;
		16'hF20F: out_word = 8'hA1;
		16'hF210: out_word = 8'hF8;
		16'hF211: out_word = 8'h1E;
		16'hF212: out_word = 8'hE0;
		16'hF213: out_word = 8'hB8;
		16'hF214: out_word = 8'h5C;
		16'hF215: out_word = 8'hE0;
		16'hF216: out_word = 8'hF0;
		16'hF217: out_word = 8'hC9;
		16'hF218: out_word = 8'h6E;
		16'hF219: out_word = 8'hF3;
		16'hF21A: out_word = 8'hE0;
		16'hF21B: out_word = 8'hC4;
		16'hF21C: out_word = 8'h40;
		16'hF21D: out_word = 8'h28;
		16'hF21E: out_word = 8'h72;
		16'hF21F: out_word = 8'h59;
		16'hF220: out_word = 8'hF6;
		16'hF221: out_word = 8'hE8;
		16'hF222: out_word = 8'h48;
		16'hF223: out_word = 8'h70;
		16'hF224: out_word = 8'h33;
		16'hF225: out_word = 8'h88;
		16'hF226: out_word = 8'hE8;
		16'hF227: out_word = 8'hD3;
		16'hF228: out_word = 8'h29;
		16'hF229: out_word = 8'hDD;
		16'hF22A: out_word = 8'h49;
		16'hF22B: out_word = 8'hF0;
		16'hF22C: out_word = 8'h6C;
		16'hF22D: out_word = 8'h18;
		16'hF22E: out_word = 8'h70;
		16'hF22F: out_word = 8'hF0;
		16'hF230: out_word = 8'h09;
		16'hF231: out_word = 8'h64;
		16'hF232: out_word = 8'hF8;
		16'hF233: out_word = 8'hB8;
		16'hF234: out_word = 8'h4C;
		16'hF235: out_word = 8'hD0;
		16'hF236: out_word = 8'h8D;
		16'hF237: out_word = 8'hCA;
		16'hF238: out_word = 8'h48;
		16'hF239: out_word = 8'hA0;
		16'hF23A: out_word = 8'hAF;
		16'hF23B: out_word = 8'hF5;
		16'hF23C: out_word = 8'hF0;
		16'hF23D: out_word = 8'h54;
		16'hF23E: out_word = 8'h7D;
		16'hF23F: out_word = 8'hA8;
		16'hF240: out_word = 8'hE2;
		16'hF241: out_word = 8'hF0;
		16'hF242: out_word = 8'hC7;
		16'hF243: out_word = 8'hE3;
		16'hF244: out_word = 8'h18;
		16'hF245: out_word = 8'h42;
		16'hF246: out_word = 8'h00;
		16'hF247: out_word = 8'hFB;
		16'hF248: out_word = 8'hBB;
		16'hF249: out_word = 8'hD7;
		16'hF24A: out_word = 8'h18;
		16'hF24B: out_word = 8'h44;
		16'hF24C: out_word = 8'h9A;
		16'hF24D: out_word = 8'hD0;
		16'hF24E: out_word = 8'h2D;
		16'hF24F: out_word = 8'hF8;
		16'hF250: out_word = 8'h28;
		16'hF251: out_word = 8'h05;
		16'hF252: out_word = 8'hF0;
		16'hF253: out_word = 8'hB7;
		16'hF254: out_word = 8'h7D;
		16'hF255: out_word = 8'h98;
		16'hF256: out_word = 8'h07;
		16'hF257: out_word = 8'hF3;
		16'hF258: out_word = 8'h05;
		16'hF259: out_word = 8'hC7;
		16'hF25A: out_word = 8'hA8;
		16'hF25B: out_word = 8'h06;
		16'hF25C: out_word = 8'hF7;
		16'hF25D: out_word = 8'h77;
		16'hF25E: out_word = 8'hF2;
		16'hF25F: out_word = 8'hE8;
		16'hF260: out_word = 8'h18;
		16'hF261: out_word = 8'h30;
		16'hF262: out_word = 8'h58;
		16'hF263: out_word = 8'h94;
		16'hF264: out_word = 8'hC0;
		16'hF265: out_word = 8'h20;
		16'hF266: out_word = 8'hFF;
		16'hF267: out_word = 8'h4D;
		16'hF268: out_word = 8'hD0;
		16'hF269: out_word = 8'h80;
		16'hF26A: out_word = 8'h40;
		16'hF26B: out_word = 8'h28;
		16'hF26C: out_word = 8'h0F;
		16'hF26D: out_word = 8'h04;
		16'hF26E: out_word = 8'hF0;
		16'hF26F: out_word = 8'hEF;
		16'hF270: out_word = 8'hA3;
		16'hF271: out_word = 8'h60;
		16'hF272: out_word = 8'hF0;
		16'hF273: out_word = 8'hCD;
		16'hF274: out_word = 8'hD3;
		16'hF275: out_word = 8'hD0;
		16'hF276: out_word = 8'hFF;
		16'hF277: out_word = 8'hFC;
		16'hF278: out_word = 8'h39;
		16'hF279: out_word = 8'h18;
		16'hF27A: out_word = 8'h24;
		16'hF27B: out_word = 8'h70;
		16'hF27C: out_word = 8'hD8;
		16'hF27D: out_word = 8'h77;
		16'hF27E: out_word = 8'hCE;
		16'hF27F: out_word = 8'hE7;
		16'hF280: out_word = 8'h91;
		16'hF281: out_word = 8'h3C;
		16'hF282: out_word = 8'h44;
		16'hF283: out_word = 8'h33;
		16'hF284: out_word = 8'h8F;
		16'hF285: out_word = 8'h50;
		16'hF286: out_word = 8'h34;
		16'hF287: out_word = 8'h00;
		16'hF288: out_word = 8'hFD;
		16'hF289: out_word = 8'hFF;
		16'hF28A: out_word = 8'h3C;
		16'hF28B: out_word = 8'h11;
		16'hF28C: out_word = 8'h30;
		16'hF28D: out_word = 8'hE9;
		16'hF28E: out_word = 8'h11;
		16'hF28F: out_word = 8'hE8;
		16'hF290: out_word = 8'hF0;
		16'hF291: out_word = 8'h00;
		16'hF292: out_word = 8'h58;
		16'hF293: out_word = 8'h72;
		16'hF294: out_word = 8'hC0;
		16'hF295: out_word = 8'h20;
		16'hF296: out_word = 8'h89;
		16'hF297: out_word = 8'hCF;
		16'hF298: out_word = 8'hF0;
		16'hF299: out_word = 8'h3C;
		16'hF29A: out_word = 8'h7F;
		16'hF29B: out_word = 8'hDC;
		16'hF29C: out_word = 8'h8F;
		16'hF29D: out_word = 8'hD0;
		16'hF29E: out_word = 8'h78;
		16'hF29F: out_word = 8'h00;
		16'hF2A0: out_word = 8'hDE;
		16'hF2A1: out_word = 8'h85;
		16'hF2A2: out_word = 8'h30;
		16'hF2A3: out_word = 8'h00;
		16'hF2A4: out_word = 8'h80;
		16'hF2A5: out_word = 8'h08;
		16'hF2A6: out_word = 8'h8B;
		16'hF2A7: out_word = 8'h98;
		16'hF2A8: out_word = 8'hD1;
		16'hF2A9: out_word = 8'h07;
		16'hF2AA: out_word = 8'h40;
		16'hF2AB: out_word = 8'h31;
		16'hF2AC: out_word = 8'h50;
		16'hF2AD: out_word = 8'h60;
		16'hF2AE: out_word = 8'h97;
		16'hF2AF: out_word = 8'h9C;
		16'hF2B0: out_word = 8'h90;
		16'hF2B1: out_word = 8'h79;
		16'hF2B2: out_word = 8'h70;
		16'hF2B3: out_word = 8'h50;
		16'hF2B4: out_word = 8'h6D;
		16'hF2B5: out_word = 8'h68;
		16'hF2B6: out_word = 8'h54;
		16'hF2B7: out_word = 8'h13;
		16'hF2B8: out_word = 8'hFF;
		16'hF2B9: out_word = 8'hF8;
		16'hF2BA: out_word = 8'h58;
		16'hF2BB: out_word = 8'h64;
		16'hF2BC: out_word = 8'h47;
		16'hF2BD: out_word = 8'hD0;
		16'hF2BE: out_word = 8'h9E;
		16'hF2BF: out_word = 8'hB0;
		16'hF2C0: out_word = 8'h30;
		16'hF2C1: out_word = 8'h6F;
		16'hF2C2: out_word = 8'hF7;
		16'hF2C3: out_word = 8'hFF;
		16'hF2C4: out_word = 8'h87;
		16'hF2C5: out_word = 8'hB0;
		16'hF2C6: out_word = 8'h71;
		16'hF2C7: out_word = 8'hE0;
		16'hF2C8: out_word = 8'hFF;
		16'hF2C9: out_word = 8'hA0;
		16'hF2CA: out_word = 8'h7F;
		16'hF2CB: out_word = 8'hD0;
		16'hF2CC: out_word = 8'hFF;
		16'hF2CD: out_word = 8'h78;
		16'hF2CE: out_word = 8'hB5;
		16'hF2CF: out_word = 8'h92;
		16'hF2D0: out_word = 8'h34;
		16'hF2D1: out_word = 8'hC0;
		16'hF2D2: out_word = 8'h3C;
		16'hF2D3: out_word = 8'h00;
		16'hF2D4: out_word = 8'h17;
		16'hF2D5: out_word = 8'hF3;
		16'hF2D6: out_word = 8'hF0;
		16'hF2D7: out_word = 8'h52;
		16'hF2D8: out_word = 8'h00;
		16'hF2D9: out_word = 8'hFB;
		16'hF2DA: out_word = 8'hFF;
		16'hF2DB: out_word = 8'h40;
		16'hF2DC: out_word = 8'h2D;
		16'hF2DD: out_word = 8'h0D;
		16'hF2DE: out_word = 8'h7D;
		16'hF2DF: out_word = 8'hFF;
		16'hF2E0: out_word = 8'h7C;
		16'hF2E1: out_word = 8'h5F;
		16'hF2E2: out_word = 8'h21;
		16'hF2E3: out_word = 8'h11;
		16'hF2E4: out_word = 8'hFE;
		16'hF2E5: out_word = 8'h68;
		16'hF2E6: out_word = 8'h8A;
		16'hF2E7: out_word = 8'h60;
		16'hF2E8: out_word = 8'hBE;
		16'hF2E9: out_word = 8'h15;
		16'hF2EA: out_word = 8'hD4;
		16'hF2EB: out_word = 8'hFF;
		16'hF2EC: out_word = 8'h4D;
		16'hF2ED: out_word = 8'hB8;
		16'hF2EE: out_word = 8'hFC;
		16'hF2EF: out_word = 8'h0C;
		16'hF2F0: out_word = 8'hDE;
		16'hF2F1: out_word = 8'hF0;
		16'hF2F2: out_word = 8'hDA;
		16'hF2F3: out_word = 8'h28;
		16'hF2F4: out_word = 8'h50;
		16'hF2F5: out_word = 8'h77;
		16'hF2F6: out_word = 8'hBD;
		16'hF2F7: out_word = 8'h84;
		16'hF2F8: out_word = 8'hB4;
		16'hF2F9: out_word = 8'h8E;
		16'hF2FA: out_word = 8'hA4;
		16'hF2FB: out_word = 8'h28;
		16'hF2FC: out_word = 8'h67;
		16'hF2FD: out_word = 8'h9F;
		16'hF2FE: out_word = 8'h1C;
		16'hF2FF: out_word = 8'h24;
		16'hF300: out_word = 8'h6B;
		16'hF301: out_word = 8'hF7;
		16'hF302: out_word = 8'h08;
		16'hF303: out_word = 8'h9B;
		16'hF304: out_word = 8'h08;
		16'hF305: out_word = 8'hFC;
		16'hF306: out_word = 8'h00;
		16'hF307: out_word = 8'hA3;
		16'hF308: out_word = 8'hB9;
		16'hF309: out_word = 8'h7A;
		16'hF30A: out_word = 8'hFF;
		16'hF30B: out_word = 8'h68;
		16'hF30C: out_word = 8'h48;
		16'hF30D: out_word = 8'h4D;
		16'hF30E: out_word = 8'hFF;
		16'hF30F: out_word = 8'hFC;
		16'hF310: out_word = 8'h84;
		16'hF311: out_word = 8'hBF;
		16'hF312: out_word = 8'hCD;
		16'hF313: out_word = 8'h00;
		16'hF314: out_word = 8'h8B;
		16'hF315: out_word = 8'h38;
		16'hF316: out_word = 8'hE3;
		16'hF317: out_word = 8'h38;
		16'hF318: out_word = 8'h41;
		16'hF319: out_word = 8'h18;
		16'hF31A: out_word = 8'h7F;
		16'hF31B: out_word = 8'hD7;
		16'hF31C: out_word = 8'h60;
		16'hF31D: out_word = 8'h64;
		16'hF31E: out_word = 8'h32;
		16'hF31F: out_word = 8'h54;
		16'hF320: out_word = 8'h2E;
		16'hF321: out_word = 8'h86;
		16'hF322: out_word = 8'h91;
		16'hF323: out_word = 8'hF3;
		16'hF324: out_word = 8'hF8;
		16'hF325: out_word = 8'h7F;
		16'hF326: out_word = 8'hA2;
		16'hF327: out_word = 8'h08;
		16'hF328: out_word = 8'hA8;
		16'hF329: out_word = 8'h00;
		16'hF32A: out_word = 8'hFF;
		16'hF32B: out_word = 8'hC9;
		16'hF32C: out_word = 8'hFB;
		16'hF32D: out_word = 8'h08;
		16'hF32E: out_word = 8'h8C;
		16'hF32F: out_word = 8'h99;
		16'hF330: out_word = 8'h9F;
		16'hF331: out_word = 8'hA2;
		16'hF332: out_word = 8'h08;
		16'hF333: out_word = 8'hF2;
		16'hF334: out_word = 8'h32;
		16'hF335: out_word = 8'hFF;
		16'hF336: out_word = 8'hBE;
		16'hF337: out_word = 8'h00;
		16'hF338: out_word = 8'h59;
		16'hF339: out_word = 8'hFA;
		16'hF33A: out_word = 8'hBF;
		16'hF33B: out_word = 8'h10;
		16'hF33C: out_word = 8'h79;
		16'hF33D: out_word = 8'h31;
		16'hF33E: out_word = 8'hC0;
		16'hF33F: out_word = 8'h92;
		16'hF340: out_word = 8'h6D;
		16'hF341: out_word = 8'h10;
		16'hF342: out_word = 8'h48;
		16'hF343: out_word = 8'h19;
		16'hF344: out_word = 8'hD0;
		16'hF345: out_word = 8'hE0;
		16'hF346: out_word = 8'h71;
		16'hF347: out_word = 8'h9B;
		16'hF348: out_word = 8'h7C;
		16'hF349: out_word = 8'h04;
		16'hF34A: out_word = 8'h40;
		16'hF34B: out_word = 8'hE0;
		16'hF34C: out_word = 8'h28;
		16'hF34D: out_word = 8'h70;
		16'hF34E: out_word = 8'hE5;
		16'hF34F: out_word = 8'hFF;
		16'hF350: out_word = 8'h7C;
		16'hF351: out_word = 8'hB0;
		16'hF352: out_word = 8'hF8;
		16'hF353: out_word = 8'hF2;
		16'hF354: out_word = 8'hEF;
		16'hF355: out_word = 8'h60;
		16'hF356: out_word = 8'h20;
		16'hF357: out_word = 8'h38;
		16'hF358: out_word = 8'h88;
		16'hF359: out_word = 8'hF6;
		16'hF35A: out_word = 8'h68;
		16'hF35B: out_word = 8'h74;
		16'hF35C: out_word = 8'h4C;
		16'hF35D: out_word = 8'h38;
		16'hF35E: out_word = 8'hAE;
		16'hF35F: out_word = 8'hF9;
		16'hF360: out_word = 8'h30;
		16'hF361: out_word = 8'h70;
		16'hF362: out_word = 8'h2E;
		16'hF363: out_word = 8'h6D;
		16'hF364: out_word = 8'h5E;
		16'hF365: out_word = 8'hA0;
		16'hF366: out_word = 8'h1C;
		16'hF367: out_word = 8'h50;
		16'hF368: out_word = 8'hE4;
		16'hF369: out_word = 8'h48;
		16'hF36A: out_word = 8'h54;
		16'hF36B: out_word = 8'h74;
		16'hF36C: out_word = 8'hD8;
		16'hF36D: out_word = 8'h36;
		16'hF36E: out_word = 8'h9F;
		16'hF36F: out_word = 8'h91;
		16'hF370: out_word = 8'h47;
		16'hF371: out_word = 8'h60;
		16'hF372: out_word = 8'hB0;
		16'hF373: out_word = 8'hF7;
		16'hF374: out_word = 8'h4C;
		16'hF375: out_word = 8'h34;
		16'hF376: out_word = 8'h2D;
		16'hF377: out_word = 8'h04;
		16'hF378: out_word = 8'hBA;
		16'hF379: out_word = 8'hA8;
		16'hF37A: out_word = 8'hFF;
		16'hF37B: out_word = 8'hBF;
		16'hF37C: out_word = 8'hFF;
		16'hF37D: out_word = 8'hE9;
		16'hF37E: out_word = 8'h00;
		16'hF37F: out_word = 8'hED;
		16'hF380: out_word = 8'h3C;
		16'hF381: out_word = 8'h2B;
		16'hF382: out_word = 8'hC1;
		16'hF383: out_word = 8'hC8;
		16'hF384: out_word = 8'hE9;
		16'hF385: out_word = 8'hE8;
		16'hF386: out_word = 8'hDF;
		16'hF387: out_word = 8'hED;
		16'hF388: out_word = 8'h00;
		16'hF389: out_word = 8'h7E;
		16'hF38A: out_word = 8'hFF;
		16'hF38B: out_word = 8'hF5;
		16'hF38C: out_word = 8'hF0;
		16'hF38D: out_word = 8'h18;
		16'hF38E: out_word = 8'hAF;
		16'hF38F: out_word = 8'hD1;
		16'hF390: out_word = 8'h70;
		16'hF391: out_word = 8'hC0;
		16'hF392: out_word = 8'h7D;
		16'hF393: out_word = 8'h91;
		16'hF394: out_word = 8'hA1;
		16'hF395: out_word = 8'hF8;
		16'hF396: out_word = 8'hAF;
		16'hF397: out_word = 8'hD2;
		16'hF398: out_word = 8'hFF;
		16'hF399: out_word = 8'hF8;
		16'hF39A: out_word = 8'h1C;
		16'hF39B: out_word = 8'hF3;
		16'hF39C: out_word = 8'h00;
		16'hF39D: out_word = 8'hFE;
		16'hF39E: out_word = 8'hFF;
		16'hF39F: out_word = 8'h8F;
		16'hF3A0: out_word = 8'h48;
		16'hF3A1: out_word = 8'hFB;
		16'hF3A2: out_word = 8'hFF;
		16'hF3A3: out_word = 8'h2F;
		16'hF3A4: out_word = 8'hF7;
		16'hF3A5: out_word = 8'h08;
		16'hF3A6: out_word = 8'h7C;
		16'hF3A7: out_word = 8'hA5;
		16'hF3A8: out_word = 8'h00;
		16'hF3A9: out_word = 8'hA8;
		16'hF3AA: out_word = 8'hB0;
		16'hF3AB: out_word = 8'hA0;
		16'hF3AC: out_word = 8'hFC;
		16'hF3AD: out_word = 8'h16;
		16'hF3AE: out_word = 8'hA8;
		16'hF3AF: out_word = 8'hFE;
		16'hF3B0: out_word = 8'hFC;
		16'hF3B1: out_word = 8'h23;
		16'hF3B2: out_word = 8'h39;
		16'hF3B3: out_word = 8'hFC;
		16'hF3B4: out_word = 8'h30;
		16'hF3B5: out_word = 8'h64;
		16'hF3B6: out_word = 8'hAD;
		16'hF3B7: out_word = 8'hFF;
		16'hF3B8: out_word = 8'hF0;
		16'hF3B9: out_word = 8'h88;
		16'hF3BA: out_word = 8'hF9;
		16'hF3BB: out_word = 8'hF7;
		16'hF3BC: out_word = 8'hED;
		16'hF3BD: out_word = 8'hC3;
		16'hF3BE: out_word = 8'hE9;
		16'hF3BF: out_word = 8'hE8;
		16'hF3C0: out_word = 8'h69;
		16'hF3C1: out_word = 8'hCB;
		16'hF3C2: out_word = 8'h5B;
		16'hF3C3: out_word = 8'hF8;
		16'hF3C4: out_word = 8'h43;
		16'hF3C5: out_word = 8'hF8;
		16'hF3C6: out_word = 8'h66;
		16'hF3C7: out_word = 8'hE8;
		16'hF3C8: out_word = 8'hE8;
		16'hF3C9: out_word = 8'h08;
		16'hF3CA: out_word = 8'h5B;
		16'hF3CB: out_word = 8'hE7;
		16'hF3CC: out_word = 8'h9C;
		16'hF3CD: out_word = 8'hFF;
		16'hF3CE: out_word = 8'hE1;
		16'hF3CF: out_word = 8'h6A;
		16'hF3D0: out_word = 8'hF0;
		16'hF3D1: out_word = 8'h32;
		16'hF3D2: out_word = 8'hE8;
		16'hF3D3: out_word = 8'hF8;
		16'hF3D4: out_word = 8'hF3;
		16'hF3D5: out_word = 8'hE0;
		16'hF3D6: out_word = 8'hF7;
		16'hF3D7: out_word = 8'h28;
		16'hF3D8: out_word = 8'hEB;
		16'hF3D9: out_word = 8'hD0;
		16'hF3DA: out_word = 8'hB8;
		16'hF3DB: out_word = 8'h8E;
		16'hF3DC: out_word = 8'hF7;
		16'hF3DD: out_word = 8'h35;
		16'hF3DE: out_word = 8'hC7;
		16'hF3DF: out_word = 8'h38;
		16'hF3E0: out_word = 8'hA0;
		16'hF3E1: out_word = 8'h2A;
		16'hF3E2: out_word = 8'hE5;
		16'hF3E3: out_word = 8'hF8;
		16'hF3E4: out_word = 8'hFC;
		16'hF3E5: out_word = 8'hB7;
		16'hF3E6: out_word = 8'h5B;
		16'hF3E7: out_word = 8'hEB;
		16'hF3E8: out_word = 8'h11;
		16'hF3E9: out_word = 8'hE8;
		16'hF3EA: out_word = 8'hFC;
		16'hF3EB: out_word = 8'hE6;
		16'hF3EC: out_word = 8'hF0;
		16'hF3ED: out_word = 8'hC6;
		16'hF3EE: out_word = 8'hE0;
		16'hF3EF: out_word = 8'hC1;
		16'hF3F0: out_word = 8'hE9;
		16'hF3F1: out_word = 8'h9A;
		16'hF3F2: out_word = 8'h2D;
		16'hF3F3: out_word = 8'h78;
		16'hF3F4: out_word = 8'h2C;
		16'hF3F5: out_word = 8'h00;
		16'hF3F6: out_word = 8'h95;
		16'hF3F7: out_word = 8'hEF;
		16'hF3F8: out_word = 8'h20;
		16'hF3F9: out_word = 8'h3C;
		16'hF3FA: out_word = 8'h04;
		16'hF3FB: out_word = 8'hC9;
		16'hF3FC: out_word = 8'h03;
		16'hF3FD: out_word = 8'h45;
		16'hF3FE: out_word = 8'hEF;
		16'hF3FF: out_word = 8'hEC;
		16'hF400: out_word = 8'h1A;
		16'hF401: out_word = 8'hCF;
		16'hF402: out_word = 8'h2D;
		16'hF403: out_word = 8'hC9;
		16'hF404: out_word = 8'hEC;
		16'hF405: out_word = 8'h48;
		16'hF406: out_word = 8'hE0;
		16'hF407: out_word = 8'hE8;
		16'hF408: out_word = 8'hF2;
		16'hF409: out_word = 8'hF0;
		16'hF40A: out_word = 8'h3C;
		16'hF40B: out_word = 8'hE8;
		16'hF40C: out_word = 8'hE0;
		16'hF40D: out_word = 8'h88;
		16'hF40E: out_word = 8'hE8;
		16'hF40F: out_word = 8'hB8;
		16'hF410: out_word = 8'hD8;
		16'hF411: out_word = 8'hF0;
		16'hF412: out_word = 8'h2B;
		16'hF413: out_word = 8'hCF;
		16'hF414: out_word = 8'hD1;
		16'hF415: out_word = 8'h35;
		16'hF416: out_word = 8'hE0;
		16'hF417: out_word = 8'h35;
		16'hF418: out_word = 8'h90;
		16'hF419: out_word = 8'h3C;
		16'hF41A: out_word = 8'h3C;
		16'hF41B: out_word = 8'h68;
		16'hF41C: out_word = 8'hF3;
		16'hF41D: out_word = 8'h90;
		16'hF41E: out_word = 8'hCF;
		16'hF41F: out_word = 8'hE0;
		16'hF420: out_word = 8'h3C;
		16'hF421: out_word = 8'h88;
		16'hF422: out_word = 8'hF7;
		16'hF423: out_word = 8'hD4;
		16'hF424: out_word = 8'hE0;
		16'hF425: out_word = 8'h8F;
		16'hF426: out_word = 8'hB9;
		16'hF427: out_word = 8'h36;
		16'hF428: out_word = 8'hB8;
		16'hF429: out_word = 8'h23;
		16'hF42A: out_word = 8'h67;
		16'hF42B: out_word = 8'h29;
		16'hF42C: out_word = 8'h52;
		16'hF42D: out_word = 8'hD7;
		16'hF42E: out_word = 8'h35;
		16'hF42F: out_word = 8'hEB;
		16'hF430: out_word = 8'h3C;
		16'hF431: out_word = 8'hFF;
		16'hF432: out_word = 8'hB0;
		16'hF433: out_word = 8'h96;
		16'hF434: out_word = 8'hFF;
		16'hF435: out_word = 8'hE0;
		16'hF436: out_word = 8'hAB;
		16'hF437: out_word = 8'hFF;
		16'hF438: out_word = 8'h1C;
		16'hF439: out_word = 8'h53;
		16'hF43A: out_word = 8'hFF;
		16'hF43B: out_word = 8'h63;
		16'hF43C: out_word = 8'hE4;
		16'hF43D: out_word = 8'h33;
		16'hF43E: out_word = 8'hC5;
		16'hF43F: out_word = 8'h7F;
		16'hF440: out_word = 8'h97;
		16'hF441: out_word = 8'hAF;
		16'hF442: out_word = 8'h91;
		16'hF443: out_word = 8'h7F;
		16'hF444: out_word = 8'hF8;
		16'hF445: out_word = 8'hB6;
		16'hF446: out_word = 8'hC4;
		16'hF447: out_word = 8'hB0;
		16'hF448: out_word = 8'h7F;
		16'hF449: out_word = 8'h9B;
		16'hF44A: out_word = 8'h80;
		16'hF44B: out_word = 8'hF5;
		16'hF44C: out_word = 8'h98;
		16'hF44D: out_word = 8'hFE;
		16'hF44E: out_word = 8'h7F;
		16'hF44F: out_word = 8'hAF;
		16'hF450: out_word = 8'h34;
		16'hF451: out_word = 8'h35;
		16'hF452: out_word = 8'h87;
		16'hF453: out_word = 8'hF0;
		16'hF454: out_word = 8'h80;
		16'hF455: out_word = 8'h0F;
		16'hF456: out_word = 8'hF3;
		16'hF457: out_word = 8'h88;
		16'hF458: out_word = 8'h62;
		16'hF459: out_word = 8'hF8;
		16'hF45A: out_word = 8'h5A;
		16'hF45B: out_word = 8'hEF;
		16'hF45C: out_word = 8'h60;
		16'hF45D: out_word = 8'h78;
		16'hF45E: out_word = 8'h80;
		16'hF45F: out_word = 8'h06;
		16'hF460: out_word = 8'hBE;
		16'hF461: out_word = 8'h80;
		16'hF462: out_word = 8'h01;
		16'hF463: out_word = 8'hAF;
		16'hF464: out_word = 8'h8C;
		16'hF465: out_word = 8'h80;
		16'hF466: out_word = 8'h98;
		16'hF467: out_word = 8'h04;
		16'hF468: out_word = 8'h88;
		16'hF469: out_word = 8'hD0;
		16'hF46A: out_word = 8'h03;
		16'hF46B: out_word = 8'h4F;
		16'hF46C: out_word = 8'h08;
		16'hF46D: out_word = 8'h7F;
		16'hF46E: out_word = 8'hE3;
		16'hF46F: out_word = 8'h5A;
		16'hF470: out_word = 8'hFD;
		16'hF471: out_word = 8'h80;
		16'hF472: out_word = 8'h28;
		16'hF473: out_word = 8'h6B;
		16'hF474: out_word = 8'hD0;
		16'hF475: out_word = 8'hA8;
		16'hF476: out_word = 8'h1A;
		16'hF477: out_word = 8'hF9;
		16'hF478: out_word = 8'hA0;
		16'hF479: out_word = 8'hFB;
		16'hF47A: out_word = 8'h61;
		16'hF47B: out_word = 8'h97;
		16'hF47C: out_word = 8'h24;
		16'hF47D: out_word = 8'hFD;
		16'hF47E: out_word = 8'hEE;
		16'hF47F: out_word = 8'h49;
		16'hF480: out_word = 8'h48;
		16'hF481: out_word = 8'h62;
		16'hF482: out_word = 8'hFD;
		16'hF483: out_word = 8'h30;
		16'hF484: out_word = 8'h3F;
		16'hF485: out_word = 8'hAB;
		16'hF486: out_word = 8'h78;
		16'hF487: out_word = 8'h8F;
		16'hF488: out_word = 8'hAB;
		16'hF489: out_word = 8'hE3;
		16'hF48A: out_word = 8'hA9;
		16'hF48B: out_word = 8'hF6;
		16'hF48C: out_word = 8'h28;
		16'hF48D: out_word = 8'h5C;
		16'hF48E: out_word = 8'hD2;
		16'hF48F: out_word = 8'h70;
		16'hF490: out_word = 8'h9D;
		16'hF491: out_word = 8'h34;
		16'hF492: out_word = 8'hBB;
		16'hF493: out_word = 8'h24;
		16'hF494: out_word = 8'h58;
		16'hF495: out_word = 8'hB6;
		16'hF496: out_word = 8'h40;
		16'hF497: out_word = 8'h89;
		16'hF498: out_word = 8'h71;
		16'hF499: out_word = 8'h57;
		16'hF49A: out_word = 8'hC6;
		16'hF49B: out_word = 8'h8A;
		16'hF49C: out_word = 8'hA7;
		16'hF49D: out_word = 8'hF5;
		16'hF49E: out_word = 8'h68;
		16'hF49F: out_word = 8'hA0;
		16'hF4A0: out_word = 8'h78;
		16'hF4A1: out_word = 8'h50;
		16'hF4A2: out_word = 8'hEB;
		16'hF4A3: out_word = 8'h88;
		16'hF4A4: out_word = 8'h58;
		16'hF4A5: out_word = 8'h82;
		16'hF4A6: out_word = 8'h88;
		16'hF4A7: out_word = 8'h92;
		16'hF4A8: out_word = 8'hD9;
		16'hF4A9: out_word = 8'h6D;
		16'hF4AA: out_word = 8'hB0;
		16'hF4AB: out_word = 8'h78;
		16'hF4AC: out_word = 8'h83;
		16'hF4AD: out_word = 8'hD8;
		16'hF4AE: out_word = 8'h3C;
		16'hF4AF: out_word = 8'h71;
		16'hF4B0: out_word = 8'h39;
		16'hF4B1: out_word = 8'hDF;
		16'hF4B2: out_word = 8'hD8;
		16'hF4B3: out_word = 8'h60;
		16'hF4B4: out_word = 8'h70;
		16'hF4B5: out_word = 8'h04;
		16'hF4B6: out_word = 8'hFF;
		16'hF4B7: out_word = 8'hFF;
		16'hF4B8: out_word = 8'hFF;
		16'hF4B9: out_word = 8'hFF;
		16'hF4BA: out_word = 8'hFF;
		16'hF4BB: out_word = 8'hFF;
		16'hF4BC: out_word = 8'hFF;
		16'hF4BD: out_word = 8'hFF;
		16'hF4BE: out_word = 8'hFF;
		16'hF4BF: out_word = 8'hFF;
		16'hF4C0: out_word = 8'hFF;
		16'hF4C1: out_word = 8'hFF;
		16'hF4C2: out_word = 8'hFF;
		16'hF4C3: out_word = 8'hFF;
		16'hF4C4: out_word = 8'hFF;
		16'hF4C5: out_word = 8'hFF;
		16'hF4C6: out_word = 8'hFF;
		16'hF4C7: out_word = 8'hFF;
		16'hF4C8: out_word = 8'hFF;
		16'hF4C9: out_word = 8'hFF;
		16'hF4CA: out_word = 8'hFF;
		16'hF4CB: out_word = 8'hFF;
		16'hF4CC: out_word = 8'hFF;
		16'hF4CD: out_word = 8'hFF;
		16'hF4CE: out_word = 8'hFF;
		16'hF4CF: out_word = 8'hFF;
		16'hF4D0: out_word = 8'hFF;
		16'hF4D1: out_word = 8'hFF;
		16'hF4D2: out_word = 8'hFF;
		16'hF4D3: out_word = 8'hFF;
		16'hF4D4: out_word = 8'hFF;
		16'hF4D5: out_word = 8'hFF;
		16'hF4D6: out_word = 8'hFF;
		16'hF4D7: out_word = 8'hFF;
		16'hF4D8: out_word = 8'hFF;
		16'hF4D9: out_word = 8'hFF;
		16'hF4DA: out_word = 8'hFF;
		16'hF4DB: out_word = 8'hFF;
		16'hF4DC: out_word = 8'hFF;
		16'hF4DD: out_word = 8'hFF;
		16'hF4DE: out_word = 8'hFF;
		16'hF4DF: out_word = 8'hFF;
		16'hF4E0: out_word = 8'hFF;
		16'hF4E1: out_word = 8'hFF;
		16'hF4E2: out_word = 8'hFF;
		16'hF4E3: out_word = 8'hFF;
		16'hF4E4: out_word = 8'hFF;
		16'hF4E5: out_word = 8'hFF;
		16'hF4E6: out_word = 8'hFF;
		16'hF4E7: out_word = 8'hFF;
		16'hF4E8: out_word = 8'hFF;
		16'hF4E9: out_word = 8'hFF;
		16'hF4EA: out_word = 8'hFF;
		16'hF4EB: out_word = 8'hFF;
		16'hF4EC: out_word = 8'hFF;
		16'hF4ED: out_word = 8'hFF;
		16'hF4EE: out_word = 8'hFF;
		16'hF4EF: out_word = 8'hFF;
		16'hF4F0: out_word = 8'hFF;
		16'hF4F1: out_word = 8'hFF;
		16'hF4F2: out_word = 8'hFF;
		16'hF4F3: out_word = 8'hFF;
		16'hF4F4: out_word = 8'hFF;
		16'hF4F5: out_word = 8'hFF;
		16'hF4F6: out_word = 8'hFF;
		16'hF4F7: out_word = 8'hFF;
		16'hF4F8: out_word = 8'hFF;
		16'hF4F9: out_word = 8'hFF;
		16'hF4FA: out_word = 8'hFF;
		16'hF4FB: out_word = 8'hFF;
		16'hF4FC: out_word = 8'hFF;
		16'hF4FD: out_word = 8'hFF;
		16'hF4FE: out_word = 8'hFF;
		16'hF4FF: out_word = 8'hFF;
		16'hF500: out_word = 8'hFF;
		16'hF501: out_word = 8'hFF;
		16'hF502: out_word = 8'hFF;
		16'hF503: out_word = 8'hFF;
		16'hF504: out_word = 8'hFF;
		16'hF505: out_word = 8'hFF;
		16'hF506: out_word = 8'hFF;
		16'hF507: out_word = 8'hFF;
		16'hF508: out_word = 8'hFF;
		16'hF509: out_word = 8'hFF;
		16'hF50A: out_word = 8'hFF;
		16'hF50B: out_word = 8'hFF;
		16'hF50C: out_word = 8'hFF;
		16'hF50D: out_word = 8'hFF;
		16'hF50E: out_word = 8'hFF;
		16'hF50F: out_word = 8'hFF;
		16'hF510: out_word = 8'hFF;
		16'hF511: out_word = 8'hFF;
		16'hF512: out_word = 8'hFF;
		16'hF513: out_word = 8'hFF;
		16'hF514: out_word = 8'hFF;
		16'hF515: out_word = 8'hFF;
		16'hF516: out_word = 8'hFF;
		16'hF517: out_word = 8'hFF;
		16'hF518: out_word = 8'hFF;
		16'hF519: out_word = 8'hFF;
		16'hF51A: out_word = 8'hFF;
		16'hF51B: out_word = 8'hFF;
		16'hF51C: out_word = 8'hFF;
		16'hF51D: out_word = 8'hFF;
		16'hF51E: out_word = 8'hFF;
		16'hF51F: out_word = 8'hFF;
		16'hF520: out_word = 8'hFF;
		16'hF521: out_word = 8'hFF;
		16'hF522: out_word = 8'hFF;
		16'hF523: out_word = 8'hFF;
		16'hF524: out_word = 8'hFF;
		16'hF525: out_word = 8'hFF;
		16'hF526: out_word = 8'hFF;
		16'hF527: out_word = 8'hFF;
		16'hF528: out_word = 8'hFF;
		16'hF529: out_word = 8'hFF;
		16'hF52A: out_word = 8'hFF;
		16'hF52B: out_word = 8'hFF;
		16'hF52C: out_word = 8'hFF;
		16'hF52D: out_word = 8'hFF;
		16'hF52E: out_word = 8'hFF;
		16'hF52F: out_word = 8'hFF;
		16'hF530: out_word = 8'hFF;
		16'hF531: out_word = 8'hFF;
		16'hF532: out_word = 8'hFF;
		16'hF533: out_word = 8'hFF;
		16'hF534: out_word = 8'hFF;
		16'hF535: out_word = 8'hFF;
		16'hF536: out_word = 8'hFF;
		16'hF537: out_word = 8'hFF;
		16'hF538: out_word = 8'hFF;
		16'hF539: out_word = 8'hFF;
		16'hF53A: out_word = 8'hFF;
		16'hF53B: out_word = 8'hFF;
		16'hF53C: out_word = 8'hFF;
		16'hF53D: out_word = 8'hFF;
		16'hF53E: out_word = 8'hFF;
		16'hF53F: out_word = 8'hFF;
		16'hF540: out_word = 8'hFF;
		16'hF541: out_word = 8'hFF;
		16'hF542: out_word = 8'hFF;
		16'hF543: out_word = 8'hFF;
		16'hF544: out_word = 8'hFF;
		16'hF545: out_word = 8'hFF;
		16'hF546: out_word = 8'hFF;
		16'hF547: out_word = 8'hFF;
		16'hF548: out_word = 8'hFF;
		16'hF549: out_word = 8'hFF;
		16'hF54A: out_word = 8'hFF;
		16'hF54B: out_word = 8'hFF;
		16'hF54C: out_word = 8'hFF;
		16'hF54D: out_word = 8'hFF;
		16'hF54E: out_word = 8'hFF;
		16'hF54F: out_word = 8'hFF;
		16'hF550: out_word = 8'hFF;
		16'hF551: out_word = 8'hFF;
		16'hF552: out_word = 8'hFF;
		16'hF553: out_word = 8'hFF;
		16'hF554: out_word = 8'hFF;
		16'hF555: out_word = 8'hFF;
		16'hF556: out_word = 8'hFF;
		16'hF557: out_word = 8'hFF;
		16'hF558: out_word = 8'hFF;
		16'hF559: out_word = 8'hFF;
		16'hF55A: out_word = 8'hFF;
		16'hF55B: out_word = 8'hFF;
		16'hF55C: out_word = 8'hFF;
		16'hF55D: out_word = 8'hFF;
		16'hF55E: out_word = 8'hFF;
		16'hF55F: out_word = 8'hFF;
		16'hF560: out_word = 8'hFF;
		16'hF561: out_word = 8'hFF;
		16'hF562: out_word = 8'hFF;
		16'hF563: out_word = 8'hFF;
		16'hF564: out_word = 8'hFF;
		16'hF565: out_word = 8'hFF;
		16'hF566: out_word = 8'hFF;
		16'hF567: out_word = 8'hFF;
		16'hF568: out_word = 8'hFF;
		16'hF569: out_word = 8'hFF;
		16'hF56A: out_word = 8'hFF;
		16'hF56B: out_word = 8'hFF;
		16'hF56C: out_word = 8'hFF;
		16'hF56D: out_word = 8'hFF;
		16'hF56E: out_word = 8'hFF;
		16'hF56F: out_word = 8'hFF;
		16'hF570: out_word = 8'hFF;
		16'hF571: out_word = 8'hFF;
		16'hF572: out_word = 8'hFF;
		16'hF573: out_word = 8'hFF;
		16'hF574: out_word = 8'hFF;
		16'hF575: out_word = 8'hFF;
		16'hF576: out_word = 8'hFF;
		16'hF577: out_word = 8'hFF;
		16'hF578: out_word = 8'hFF;
		16'hF579: out_word = 8'hFF;
		16'hF57A: out_word = 8'hFF;
		16'hF57B: out_word = 8'hFF;
		16'hF57C: out_word = 8'hFF;
		16'hF57D: out_word = 8'hFF;
		16'hF57E: out_word = 8'hFF;
		16'hF57F: out_word = 8'hFF;
		16'hF580: out_word = 8'hFF;
		16'hF581: out_word = 8'hFF;
		16'hF582: out_word = 8'hFF;
		16'hF583: out_word = 8'hFF;
		16'hF584: out_word = 8'hFF;
		16'hF585: out_word = 8'hFF;
		16'hF586: out_word = 8'hFF;
		16'hF587: out_word = 8'hFF;
		16'hF588: out_word = 8'hFF;
		16'hF589: out_word = 8'hFF;
		16'hF58A: out_word = 8'hFF;
		16'hF58B: out_word = 8'hFF;
		16'hF58C: out_word = 8'hFF;
		16'hF58D: out_word = 8'hFF;
		16'hF58E: out_word = 8'hFF;
		16'hF58F: out_word = 8'hFF;
		16'hF590: out_word = 8'hFF;
		16'hF591: out_word = 8'hFF;
		16'hF592: out_word = 8'hFF;
		16'hF593: out_word = 8'hFF;
		16'hF594: out_word = 8'hFF;
		16'hF595: out_word = 8'hFF;
		16'hF596: out_word = 8'hFF;
		16'hF597: out_word = 8'hFF;
		16'hF598: out_word = 8'hFF;
		16'hF599: out_word = 8'hFF;
		16'hF59A: out_word = 8'hFF;
		16'hF59B: out_word = 8'hFF;
		16'hF59C: out_word = 8'hFF;
		16'hF59D: out_word = 8'hFF;
		16'hF59E: out_word = 8'hFF;
		16'hF59F: out_word = 8'hFF;
		16'hF5A0: out_word = 8'hFF;
		16'hF5A1: out_word = 8'hFF;
		16'hF5A2: out_word = 8'hFF;
		16'hF5A3: out_word = 8'hFF;
		16'hF5A4: out_word = 8'hFF;
		16'hF5A5: out_word = 8'hFF;
		16'hF5A6: out_word = 8'hFF;
		16'hF5A7: out_word = 8'hFF;
		16'hF5A8: out_word = 8'hFF;
		16'hF5A9: out_word = 8'hFF;
		16'hF5AA: out_word = 8'hFF;
		16'hF5AB: out_word = 8'hFF;
		16'hF5AC: out_word = 8'hFF;
		16'hF5AD: out_word = 8'hFF;
		16'hF5AE: out_word = 8'hFF;
		16'hF5AF: out_word = 8'hFF;
		16'hF5B0: out_word = 8'hFF;
		16'hF5B1: out_word = 8'hFF;
		16'hF5B2: out_word = 8'hFF;
		16'hF5B3: out_word = 8'hFF;
		16'hF5B4: out_word = 8'hFF;
		16'hF5B5: out_word = 8'hFF;
		16'hF5B6: out_word = 8'hFF;
		16'hF5B7: out_word = 8'hFF;
		16'hF5B8: out_word = 8'hFF;
		16'hF5B9: out_word = 8'hFF;
		16'hF5BA: out_word = 8'hFF;
		16'hF5BB: out_word = 8'hFF;
		16'hF5BC: out_word = 8'hFF;
		16'hF5BD: out_word = 8'hFF;
		16'hF5BE: out_word = 8'hFF;
		16'hF5BF: out_word = 8'hFF;
		16'hF5C0: out_word = 8'hFF;
		16'hF5C1: out_word = 8'hFF;
		16'hF5C2: out_word = 8'hFF;
		16'hF5C3: out_word = 8'hFF;
		16'hF5C4: out_word = 8'hFF;
		16'hF5C5: out_word = 8'hFF;
		16'hF5C6: out_word = 8'hFF;
		16'hF5C7: out_word = 8'hFF;
		16'hF5C8: out_word = 8'hFF;
		16'hF5C9: out_word = 8'hFF;
		16'hF5CA: out_word = 8'hFF;
		16'hF5CB: out_word = 8'hFF;
		16'hF5CC: out_word = 8'hFF;
		16'hF5CD: out_word = 8'hFF;
		16'hF5CE: out_word = 8'hFF;
		16'hF5CF: out_word = 8'hFF;
		16'hF5D0: out_word = 8'hFF;
		16'hF5D1: out_word = 8'hFF;
		16'hF5D2: out_word = 8'hFF;
		16'hF5D3: out_word = 8'hFF;
		16'hF5D4: out_word = 8'hFF;
		16'hF5D5: out_word = 8'hFF;
		16'hF5D6: out_word = 8'hFF;
		16'hF5D7: out_word = 8'hFF;
		16'hF5D8: out_word = 8'hFF;
		16'hF5D9: out_word = 8'hFF;
		16'hF5DA: out_word = 8'hFF;
		16'hF5DB: out_word = 8'hFF;
		16'hF5DC: out_word = 8'hFF;
		16'hF5DD: out_word = 8'hFF;
		16'hF5DE: out_word = 8'hFF;
		16'hF5DF: out_word = 8'hFF;
		16'hF5E0: out_word = 8'hFF;
		16'hF5E1: out_word = 8'hFF;
		16'hF5E2: out_word = 8'hFF;
		16'hF5E3: out_word = 8'hFF;
		16'hF5E4: out_word = 8'hFF;
		16'hF5E5: out_word = 8'hFF;
		16'hF5E6: out_word = 8'hFF;
		16'hF5E7: out_word = 8'hFF;
		16'hF5E8: out_word = 8'hFF;
		16'hF5E9: out_word = 8'hFF;
		16'hF5EA: out_word = 8'hFF;
		16'hF5EB: out_word = 8'hFF;
		16'hF5EC: out_word = 8'hFF;
		16'hF5ED: out_word = 8'hFF;
		16'hF5EE: out_word = 8'hFF;
		16'hF5EF: out_word = 8'hFF;
		16'hF5F0: out_word = 8'hFF;
		16'hF5F1: out_word = 8'hFF;
		16'hF5F2: out_word = 8'hFF;
		16'hF5F3: out_word = 8'hFF;
		16'hF5F4: out_word = 8'hFF;
		16'hF5F5: out_word = 8'hFF;
		16'hF5F6: out_word = 8'hFF;
		16'hF5F7: out_word = 8'hFF;
		16'hF5F8: out_word = 8'hFF;
		16'hF5F9: out_word = 8'hFF;
		16'hF5FA: out_word = 8'hFF;
		16'hF5FB: out_word = 8'hFF;
		16'hF5FC: out_word = 8'hFF;
		16'hF5FD: out_word = 8'hFF;
		16'hF5FE: out_word = 8'hFF;
		16'hF5FF: out_word = 8'hFF;
		16'hF600: out_word = 8'hFF;
		16'hF601: out_word = 8'hFF;
		16'hF602: out_word = 8'hFF;
		16'hF603: out_word = 8'hFF;
		16'hF604: out_word = 8'hFF;
		16'hF605: out_word = 8'hFF;
		16'hF606: out_word = 8'hFF;
		16'hF607: out_word = 8'hFF;
		16'hF608: out_word = 8'hFF;
		16'hF609: out_word = 8'hFF;
		16'hF60A: out_word = 8'hFF;
		16'hF60B: out_word = 8'hFF;
		16'hF60C: out_word = 8'hFF;
		16'hF60D: out_word = 8'hFF;
		16'hF60E: out_word = 8'hFF;
		16'hF60F: out_word = 8'hFF;
		16'hF610: out_word = 8'hFF;
		16'hF611: out_word = 8'hFF;
		16'hF612: out_word = 8'hFF;
		16'hF613: out_word = 8'hFF;
		16'hF614: out_word = 8'hFF;
		16'hF615: out_word = 8'hFF;
		16'hF616: out_word = 8'hFF;
		16'hF617: out_word = 8'hFF;
		16'hF618: out_word = 8'hFF;
		16'hF619: out_word = 8'hFF;
		16'hF61A: out_word = 8'hFF;
		16'hF61B: out_word = 8'hFF;
		16'hF61C: out_word = 8'hFF;
		16'hF61D: out_word = 8'hFF;
		16'hF61E: out_word = 8'hFF;
		16'hF61F: out_word = 8'hFF;
		16'hF620: out_word = 8'hFF;
		16'hF621: out_word = 8'hFF;
		16'hF622: out_word = 8'hFF;
		16'hF623: out_word = 8'hFF;
		16'hF624: out_word = 8'hFF;
		16'hF625: out_word = 8'hFF;
		16'hF626: out_word = 8'hFF;
		16'hF627: out_word = 8'hFF;
		16'hF628: out_word = 8'hFF;
		16'hF629: out_word = 8'hFF;
		16'hF62A: out_word = 8'hFF;
		16'hF62B: out_word = 8'hFF;
		16'hF62C: out_word = 8'hFF;
		16'hF62D: out_word = 8'hFF;
		16'hF62E: out_word = 8'hFF;
		16'hF62F: out_word = 8'hFF;
		16'hF630: out_word = 8'hFF;
		16'hF631: out_word = 8'hFF;
		16'hF632: out_word = 8'hFF;
		16'hF633: out_word = 8'hFF;
		16'hF634: out_word = 8'hFF;
		16'hF635: out_word = 8'hFF;
		16'hF636: out_word = 8'hFF;
		16'hF637: out_word = 8'hFF;
		16'hF638: out_word = 8'hFF;
		16'hF639: out_word = 8'hFF;
		16'hF63A: out_word = 8'hFF;
		16'hF63B: out_word = 8'hFF;
		16'hF63C: out_word = 8'hFF;
		16'hF63D: out_word = 8'hFF;
		16'hF63E: out_word = 8'hFF;
		16'hF63F: out_word = 8'hFF;
		16'hF640: out_word = 8'hFF;
		16'hF641: out_word = 8'hFF;
		16'hF642: out_word = 8'hFF;
		16'hF643: out_word = 8'hFF;
		16'hF644: out_word = 8'hFF;
		16'hF645: out_word = 8'hFF;
		16'hF646: out_word = 8'hFF;
		16'hF647: out_word = 8'hFF;
		16'hF648: out_word = 8'hFF;
		16'hF649: out_word = 8'hFF;
		16'hF64A: out_word = 8'hFF;
		16'hF64B: out_word = 8'hFF;
		16'hF64C: out_word = 8'hFF;
		16'hF64D: out_word = 8'hFF;
		16'hF64E: out_word = 8'hFF;
		16'hF64F: out_word = 8'hFF;
		16'hF650: out_word = 8'hFF;
		16'hF651: out_word = 8'hFF;
		16'hF652: out_word = 8'hFF;
		16'hF653: out_word = 8'hFF;
		16'hF654: out_word = 8'hFF;
		16'hF655: out_word = 8'hFF;
		16'hF656: out_word = 8'hFF;
		16'hF657: out_word = 8'hFF;
		16'hF658: out_word = 8'hFF;
		16'hF659: out_word = 8'hFF;
		16'hF65A: out_word = 8'hFF;
		16'hF65B: out_word = 8'hFF;
		16'hF65C: out_word = 8'hFF;
		16'hF65D: out_word = 8'hFF;
		16'hF65E: out_word = 8'hFF;
		16'hF65F: out_word = 8'hFF;
		16'hF660: out_word = 8'hFF;
		16'hF661: out_word = 8'hFF;
		16'hF662: out_word = 8'hFF;
		16'hF663: out_word = 8'hFF;
		16'hF664: out_word = 8'hFF;
		16'hF665: out_word = 8'hFF;
		16'hF666: out_word = 8'hFF;
		16'hF667: out_word = 8'hFF;
		16'hF668: out_word = 8'hFF;
		16'hF669: out_word = 8'hFF;
		16'hF66A: out_word = 8'hFF;
		16'hF66B: out_word = 8'hFF;
		16'hF66C: out_word = 8'hFF;
		16'hF66D: out_word = 8'hFF;
		16'hF66E: out_word = 8'hFF;
		16'hF66F: out_word = 8'hFF;
		16'hF670: out_word = 8'hFF;
		16'hF671: out_word = 8'hFF;
		16'hF672: out_word = 8'hFF;
		16'hF673: out_word = 8'hFF;
		16'hF674: out_word = 8'hFF;
		16'hF675: out_word = 8'hFF;
		16'hF676: out_word = 8'hFF;
		16'hF677: out_word = 8'hFF;
		16'hF678: out_word = 8'hFF;
		16'hF679: out_word = 8'hFF;
		16'hF67A: out_word = 8'hFF;
		16'hF67B: out_word = 8'hFF;
		16'hF67C: out_word = 8'hFF;
		16'hF67D: out_word = 8'hFF;
		16'hF67E: out_word = 8'hFF;
		16'hF67F: out_word = 8'hFF;
		16'hF680: out_word = 8'hFF;
		16'hF681: out_word = 8'hFF;
		16'hF682: out_word = 8'hFF;
		16'hF683: out_word = 8'hFF;
		16'hF684: out_word = 8'hFF;
		16'hF685: out_word = 8'hFF;
		16'hF686: out_word = 8'hFF;
		16'hF687: out_word = 8'hFF;
		16'hF688: out_word = 8'hFF;
		16'hF689: out_word = 8'hFF;
		16'hF68A: out_word = 8'hFF;
		16'hF68B: out_word = 8'hFF;
		16'hF68C: out_word = 8'hFF;
		16'hF68D: out_word = 8'hFF;
		16'hF68E: out_word = 8'hFF;
		16'hF68F: out_word = 8'hFF;
		16'hF690: out_word = 8'hFF;
		16'hF691: out_word = 8'hFF;
		16'hF692: out_word = 8'hFF;
		16'hF693: out_word = 8'hFF;
		16'hF694: out_word = 8'hFF;
		16'hF695: out_word = 8'hFF;
		16'hF696: out_word = 8'hFF;
		16'hF697: out_word = 8'hFF;
		16'hF698: out_word = 8'hFF;
		16'hF699: out_word = 8'hFF;
		16'hF69A: out_word = 8'hFF;
		16'hF69B: out_word = 8'hFF;
		16'hF69C: out_word = 8'hFF;
		16'hF69D: out_word = 8'hFF;
		16'hF69E: out_word = 8'hFF;
		16'hF69F: out_word = 8'hFF;
		16'hF6A0: out_word = 8'hFF;
		16'hF6A1: out_word = 8'hFF;
		16'hF6A2: out_word = 8'hFF;
		16'hF6A3: out_word = 8'hFF;
		16'hF6A4: out_word = 8'hFF;
		16'hF6A5: out_word = 8'hFF;
		16'hF6A6: out_word = 8'hFF;
		16'hF6A7: out_word = 8'hFF;
		16'hF6A8: out_word = 8'hFF;
		16'hF6A9: out_word = 8'hFF;
		16'hF6AA: out_word = 8'hFF;
		16'hF6AB: out_word = 8'hFF;
		16'hF6AC: out_word = 8'hFF;
		16'hF6AD: out_word = 8'hFF;
		16'hF6AE: out_word = 8'hFF;
		16'hF6AF: out_word = 8'hFF;
		16'hF6B0: out_word = 8'hFF;
		16'hF6B1: out_word = 8'hFF;
		16'hF6B2: out_word = 8'hFF;
		16'hF6B3: out_word = 8'hFF;
		16'hF6B4: out_word = 8'hFF;
		16'hF6B5: out_word = 8'hFF;
		16'hF6B6: out_word = 8'hFF;
		16'hF6B7: out_word = 8'hFF;
		16'hF6B8: out_word = 8'hFF;
		16'hF6B9: out_word = 8'hFF;
		16'hF6BA: out_word = 8'hFF;
		16'hF6BB: out_word = 8'hFF;
		16'hF6BC: out_word = 8'hFF;
		16'hF6BD: out_word = 8'hFF;
		16'hF6BE: out_word = 8'hFF;
		16'hF6BF: out_word = 8'hFF;
		16'hF6C0: out_word = 8'hFF;
		16'hF6C1: out_word = 8'hFF;
		16'hF6C2: out_word = 8'hFF;
		16'hF6C3: out_word = 8'hFF;
		16'hF6C4: out_word = 8'hFF;
		16'hF6C5: out_word = 8'hFF;
		16'hF6C6: out_word = 8'hFF;
		16'hF6C7: out_word = 8'hFF;
		16'hF6C8: out_word = 8'hFF;
		16'hF6C9: out_word = 8'hFF;
		16'hF6CA: out_word = 8'hFF;
		16'hF6CB: out_word = 8'hFF;
		16'hF6CC: out_word = 8'hFF;
		16'hF6CD: out_word = 8'hFF;
		16'hF6CE: out_word = 8'hFF;
		16'hF6CF: out_word = 8'hFF;
		16'hF6D0: out_word = 8'hFF;
		16'hF6D1: out_word = 8'hFF;
		16'hF6D2: out_word = 8'hFF;
		16'hF6D3: out_word = 8'hFF;
		16'hF6D4: out_word = 8'hFF;
		16'hF6D5: out_word = 8'hFF;
		16'hF6D6: out_word = 8'hFF;
		16'hF6D7: out_word = 8'hFF;
		16'hF6D8: out_word = 8'hFF;
		16'hF6D9: out_word = 8'hFF;
		16'hF6DA: out_word = 8'hFF;
		16'hF6DB: out_word = 8'hFF;
		16'hF6DC: out_word = 8'hFF;
		16'hF6DD: out_word = 8'hFF;
		16'hF6DE: out_word = 8'hFF;
		16'hF6DF: out_word = 8'hFF;
		16'hF6E0: out_word = 8'hFF;
		16'hF6E1: out_word = 8'hFF;
		16'hF6E2: out_word = 8'hFF;
		16'hF6E3: out_word = 8'hFF;
		16'hF6E4: out_word = 8'hFF;
		16'hF6E5: out_word = 8'hFF;
		16'hF6E6: out_word = 8'hFF;
		16'hF6E7: out_word = 8'hFF;
		16'hF6E8: out_word = 8'hFF;
		16'hF6E9: out_word = 8'hFF;
		16'hF6EA: out_word = 8'hFF;
		16'hF6EB: out_word = 8'hFF;
		16'hF6EC: out_word = 8'hFF;
		16'hF6ED: out_word = 8'hFF;
		16'hF6EE: out_word = 8'hFF;
		16'hF6EF: out_word = 8'hFF;
		16'hF6F0: out_word = 8'hFF;
		16'hF6F1: out_word = 8'hFF;
		16'hF6F2: out_word = 8'hFF;
		16'hF6F3: out_word = 8'hFF;
		16'hF6F4: out_word = 8'hFF;
		16'hF6F5: out_word = 8'hFF;
		16'hF6F6: out_word = 8'hFF;
		16'hF6F7: out_word = 8'hFF;
		16'hF6F8: out_word = 8'hFF;
		16'hF6F9: out_word = 8'hFF;
		16'hF6FA: out_word = 8'hFF;
		16'hF6FB: out_word = 8'hFF;
		16'hF6FC: out_word = 8'hFF;
		16'hF6FD: out_word = 8'hFF;
		16'hF6FE: out_word = 8'hFF;
		16'hF6FF: out_word = 8'hFF;
		16'hF700: out_word = 8'hFF;
		16'hF701: out_word = 8'hFF;
		16'hF702: out_word = 8'hFF;
		16'hF703: out_word = 8'hFF;
		16'hF704: out_word = 8'hFF;
		16'hF705: out_word = 8'hFF;
		16'hF706: out_word = 8'hFF;
		16'hF707: out_word = 8'hFF;
		16'hF708: out_word = 8'hFF;
		16'hF709: out_word = 8'hFF;
		16'hF70A: out_word = 8'hFF;
		16'hF70B: out_word = 8'hFF;
		16'hF70C: out_word = 8'hFF;
		16'hF70D: out_word = 8'hFF;
		16'hF70E: out_word = 8'hFF;
		16'hF70F: out_word = 8'hFF;
		16'hF710: out_word = 8'hFF;
		16'hF711: out_word = 8'hFF;
		16'hF712: out_word = 8'hFF;
		16'hF713: out_word = 8'hFF;
		16'hF714: out_word = 8'hFF;
		16'hF715: out_word = 8'hFF;
		16'hF716: out_word = 8'hFF;
		16'hF717: out_word = 8'hFF;
		16'hF718: out_word = 8'hFF;
		16'hF719: out_word = 8'hFF;
		16'hF71A: out_word = 8'hFF;
		16'hF71B: out_word = 8'hFF;
		16'hF71C: out_word = 8'hFF;
		16'hF71D: out_word = 8'hFF;
		16'hF71E: out_word = 8'hFF;
		16'hF71F: out_word = 8'hFF;
		16'hF720: out_word = 8'hFF;
		16'hF721: out_word = 8'hFF;
		16'hF722: out_word = 8'hFF;
		16'hF723: out_word = 8'hFF;
		16'hF724: out_word = 8'hFF;
		16'hF725: out_word = 8'hFF;
		16'hF726: out_word = 8'hFF;
		16'hF727: out_word = 8'hFF;
		16'hF728: out_word = 8'hFF;
		16'hF729: out_word = 8'hFF;
		16'hF72A: out_word = 8'hFF;
		16'hF72B: out_word = 8'hFF;
		16'hF72C: out_word = 8'hFF;
		16'hF72D: out_word = 8'hFF;
		16'hF72E: out_word = 8'hFF;
		16'hF72F: out_word = 8'hFF;
		16'hF730: out_word = 8'hFF;
		16'hF731: out_word = 8'hFF;
		16'hF732: out_word = 8'hFF;
		16'hF733: out_word = 8'hFF;
		16'hF734: out_word = 8'hFF;
		16'hF735: out_word = 8'hFF;
		16'hF736: out_word = 8'hFF;
		16'hF737: out_word = 8'hFF;
		16'hF738: out_word = 8'hFF;
		16'hF739: out_word = 8'hFF;
		16'hF73A: out_word = 8'hFF;
		16'hF73B: out_word = 8'hFF;
		16'hF73C: out_word = 8'hFF;
		16'hF73D: out_word = 8'hFF;
		16'hF73E: out_word = 8'hFF;
		16'hF73F: out_word = 8'hFF;
		16'hF740: out_word = 8'hFF;
		16'hF741: out_word = 8'hFF;
		16'hF742: out_word = 8'hFF;
		16'hF743: out_word = 8'hFF;
		16'hF744: out_word = 8'hFF;
		16'hF745: out_word = 8'hFF;
		16'hF746: out_word = 8'hFF;
		16'hF747: out_word = 8'hFF;
		16'hF748: out_word = 8'hFF;
		16'hF749: out_word = 8'hFF;
		16'hF74A: out_word = 8'hFF;
		16'hF74B: out_word = 8'hFF;
		16'hF74C: out_word = 8'hFF;
		16'hF74D: out_word = 8'hFF;
		16'hF74E: out_word = 8'hFF;
		16'hF74F: out_word = 8'hFF;
		16'hF750: out_word = 8'hFF;
		16'hF751: out_word = 8'hFF;
		16'hF752: out_word = 8'hFF;
		16'hF753: out_word = 8'hFF;
		16'hF754: out_word = 8'hFF;
		16'hF755: out_word = 8'hFF;
		16'hF756: out_word = 8'hFF;
		16'hF757: out_word = 8'hFF;
		16'hF758: out_word = 8'hFF;
		16'hF759: out_word = 8'hFF;
		16'hF75A: out_word = 8'hFF;
		16'hF75B: out_word = 8'hFF;
		16'hF75C: out_word = 8'hFF;
		16'hF75D: out_word = 8'hFF;
		16'hF75E: out_word = 8'hFF;
		16'hF75F: out_word = 8'hFF;
		16'hF760: out_word = 8'hFF;
		16'hF761: out_word = 8'hFF;
		16'hF762: out_word = 8'hFF;
		16'hF763: out_word = 8'hFF;
		16'hF764: out_word = 8'hFF;
		16'hF765: out_word = 8'hFF;
		16'hF766: out_word = 8'hFF;
		16'hF767: out_word = 8'hFF;
		16'hF768: out_word = 8'hFF;
		16'hF769: out_word = 8'hFF;
		16'hF76A: out_word = 8'hFF;
		16'hF76B: out_word = 8'hFF;
		16'hF76C: out_word = 8'hFF;
		16'hF76D: out_word = 8'hFF;
		16'hF76E: out_word = 8'hFF;
		16'hF76F: out_word = 8'hFF;
		16'hF770: out_word = 8'hFF;
		16'hF771: out_word = 8'hFF;
		16'hF772: out_word = 8'hFF;
		16'hF773: out_word = 8'hFF;
		16'hF774: out_word = 8'hFF;
		16'hF775: out_word = 8'hFF;
		16'hF776: out_word = 8'hFF;
		16'hF777: out_word = 8'hFF;
		16'hF778: out_word = 8'hFF;
		16'hF779: out_word = 8'hFF;
		16'hF77A: out_word = 8'hFF;
		16'hF77B: out_word = 8'hFF;
		16'hF77C: out_word = 8'hFF;
		16'hF77D: out_word = 8'hFF;
		16'hF77E: out_word = 8'hFF;
		16'hF77F: out_word = 8'hFF;
		16'hF780: out_word = 8'hFF;
		16'hF781: out_word = 8'hFF;
		16'hF782: out_word = 8'hFF;
		16'hF783: out_word = 8'hFF;
		16'hF784: out_word = 8'hFF;
		16'hF785: out_word = 8'hFF;
		16'hF786: out_word = 8'hFF;
		16'hF787: out_word = 8'hFF;
		16'hF788: out_word = 8'hFF;
		16'hF789: out_word = 8'hFF;
		16'hF78A: out_word = 8'hFF;
		16'hF78B: out_word = 8'hFF;
		16'hF78C: out_word = 8'hFF;
		16'hF78D: out_word = 8'hFF;
		16'hF78E: out_word = 8'hFF;
		16'hF78F: out_word = 8'hFF;
		16'hF790: out_word = 8'hFF;
		16'hF791: out_word = 8'hFF;
		16'hF792: out_word = 8'hFF;
		16'hF793: out_word = 8'hFF;
		16'hF794: out_word = 8'hFF;
		16'hF795: out_word = 8'hFF;
		16'hF796: out_word = 8'hFF;
		16'hF797: out_word = 8'hFF;
		16'hF798: out_word = 8'hFF;
		16'hF799: out_word = 8'hFF;
		16'hF79A: out_word = 8'hFF;
		16'hF79B: out_word = 8'hFF;
		16'hF79C: out_word = 8'hFF;
		16'hF79D: out_word = 8'hFF;
		16'hF79E: out_word = 8'hFF;
		16'hF79F: out_word = 8'hFF;
		16'hF7A0: out_word = 8'hFF;
		16'hF7A1: out_word = 8'hFF;
		16'hF7A2: out_word = 8'hFF;
		16'hF7A3: out_word = 8'hFF;
		16'hF7A4: out_word = 8'hFF;
		16'hF7A5: out_word = 8'hFF;
		16'hF7A6: out_word = 8'hFF;
		16'hF7A7: out_word = 8'hFF;
		16'hF7A8: out_word = 8'hFF;
		16'hF7A9: out_word = 8'hFF;
		16'hF7AA: out_word = 8'hFF;
		16'hF7AB: out_word = 8'hFF;
		16'hF7AC: out_word = 8'hFF;
		16'hF7AD: out_word = 8'hFF;
		16'hF7AE: out_word = 8'hFF;
		16'hF7AF: out_word = 8'hFF;
		16'hF7B0: out_word = 8'hFF;
		16'hF7B1: out_word = 8'hFF;
		16'hF7B2: out_word = 8'hFF;
		16'hF7B3: out_word = 8'hFF;
		16'hF7B4: out_word = 8'hFF;
		16'hF7B5: out_word = 8'hFF;
		16'hF7B6: out_word = 8'hFF;
		16'hF7B7: out_word = 8'hFF;
		16'hF7B8: out_word = 8'hFF;
		16'hF7B9: out_word = 8'hFF;
		16'hF7BA: out_word = 8'hFF;
		16'hF7BB: out_word = 8'hFF;
		16'hF7BC: out_word = 8'hFF;
		16'hF7BD: out_word = 8'hFF;
		16'hF7BE: out_word = 8'hFF;
		16'hF7BF: out_word = 8'hFF;
		16'hF7C0: out_word = 8'hFF;
		16'hF7C1: out_word = 8'hFF;
		16'hF7C2: out_word = 8'hFF;
		16'hF7C3: out_word = 8'hFF;
		16'hF7C4: out_word = 8'hFF;
		16'hF7C5: out_word = 8'hFF;
		16'hF7C6: out_word = 8'hFF;
		16'hF7C7: out_word = 8'hFF;
		16'hF7C8: out_word = 8'hFF;
		16'hF7C9: out_word = 8'hFF;
		16'hF7CA: out_word = 8'hFF;
		16'hF7CB: out_word = 8'hFF;
		16'hF7CC: out_word = 8'hFF;
		16'hF7CD: out_word = 8'hFF;
		16'hF7CE: out_word = 8'hFF;
		16'hF7CF: out_word = 8'hFF;
		16'hF7D0: out_word = 8'hFF;
		16'hF7D1: out_word = 8'hFF;
		16'hF7D2: out_word = 8'hFF;
		16'hF7D3: out_word = 8'hFF;
		16'hF7D4: out_word = 8'hFF;
		16'hF7D5: out_word = 8'hFF;
		16'hF7D6: out_word = 8'hFF;
		16'hF7D7: out_word = 8'hFF;
		16'hF7D8: out_word = 8'hFF;
		16'hF7D9: out_word = 8'hFF;
		16'hF7DA: out_word = 8'hFF;
		16'hF7DB: out_word = 8'hFF;
		16'hF7DC: out_word = 8'hFF;
		16'hF7DD: out_word = 8'hFF;
		16'hF7DE: out_word = 8'hFF;
		16'hF7DF: out_word = 8'hFF;
		16'hF7E0: out_word = 8'hFF;
		16'hF7E1: out_word = 8'hFF;
		16'hF7E2: out_word = 8'hFF;
		16'hF7E3: out_word = 8'hFF;
		16'hF7E4: out_word = 8'hFF;
		16'hF7E5: out_word = 8'hFF;
		16'hF7E6: out_word = 8'hFF;
		16'hF7E7: out_word = 8'hFF;
		16'hF7E8: out_word = 8'hFF;
		16'hF7E9: out_word = 8'hFF;
		16'hF7EA: out_word = 8'hFF;
		16'hF7EB: out_word = 8'hFF;
		16'hF7EC: out_word = 8'hFF;
		16'hF7ED: out_word = 8'hFF;
		16'hF7EE: out_word = 8'hFF;
		16'hF7EF: out_word = 8'hFF;
		16'hF7F0: out_word = 8'hFF;
		16'hF7F1: out_word = 8'hFF;
		16'hF7F2: out_word = 8'hFF;
		16'hF7F3: out_word = 8'hFF;
		16'hF7F4: out_word = 8'hFF;
		16'hF7F5: out_word = 8'hFF;
		16'hF7F6: out_word = 8'hFF;
		16'hF7F7: out_word = 8'hFF;
		16'hF7F8: out_word = 8'hFF;
		16'hF7F9: out_word = 8'hFF;
		16'hF7FA: out_word = 8'hFF;
		16'hF7FB: out_word = 8'hFF;
		16'hF7FC: out_word = 8'hFF;
		16'hF7FD: out_word = 8'hFF;
		16'hF7FE: out_word = 8'hFF;
		16'hF7FF: out_word = 8'hFF;
		16'hF800: out_word = 8'hFF;
		16'hF801: out_word = 8'hFF;
		16'hF802: out_word = 8'hFF;
		16'hF803: out_word = 8'hFF;
		16'hF804: out_word = 8'hFF;
		16'hF805: out_word = 8'hFF;
		16'hF806: out_word = 8'hFF;
		16'hF807: out_word = 8'hFF;
		16'hF808: out_word = 8'hFF;
		16'hF809: out_word = 8'hFF;
		16'hF80A: out_word = 8'hFF;
		16'hF80B: out_word = 8'hFF;
		16'hF80C: out_word = 8'hFF;
		16'hF80D: out_word = 8'hFF;
		16'hF80E: out_word = 8'hFF;
		16'hF80F: out_word = 8'hFF;
		16'hF810: out_word = 8'hFF;
		16'hF811: out_word = 8'hFF;
		16'hF812: out_word = 8'hFF;
		16'hF813: out_word = 8'hFF;
		16'hF814: out_word = 8'hFF;
		16'hF815: out_word = 8'hFF;
		16'hF816: out_word = 8'hFF;
		16'hF817: out_word = 8'hFF;
		16'hF818: out_word = 8'hFF;
		16'hF819: out_word = 8'hFF;
		16'hF81A: out_word = 8'hFF;
		16'hF81B: out_word = 8'hFF;
		16'hF81C: out_word = 8'hFF;
		16'hF81D: out_word = 8'hFF;
		16'hF81E: out_word = 8'hFF;
		16'hF81F: out_word = 8'hFF;
		16'hF820: out_word = 8'hFF;
		16'hF821: out_word = 8'hFF;
		16'hF822: out_word = 8'hFF;
		16'hF823: out_word = 8'hFF;
		16'hF824: out_word = 8'hFF;
		16'hF825: out_word = 8'hFF;
		16'hF826: out_word = 8'hFF;
		16'hF827: out_word = 8'hFF;
		16'hF828: out_word = 8'hFF;
		16'hF829: out_word = 8'hFF;
		16'hF82A: out_word = 8'hFF;
		16'hF82B: out_word = 8'hFF;
		16'hF82C: out_word = 8'hFF;
		16'hF82D: out_word = 8'hFF;
		16'hF82E: out_word = 8'hFF;
		16'hF82F: out_word = 8'hFF;
		16'hF830: out_word = 8'hFF;
		16'hF831: out_word = 8'hFF;
		16'hF832: out_word = 8'hFF;
		16'hF833: out_word = 8'hFF;
		16'hF834: out_word = 8'hFF;
		16'hF835: out_word = 8'hFF;
		16'hF836: out_word = 8'hFF;
		16'hF837: out_word = 8'hFF;
		16'hF838: out_word = 8'hFF;
		16'hF839: out_word = 8'hFF;
		16'hF83A: out_word = 8'hFF;
		16'hF83B: out_word = 8'hFF;
		16'hF83C: out_word = 8'hFF;
		16'hF83D: out_word = 8'hFF;
		16'hF83E: out_word = 8'hFF;
		16'hF83F: out_word = 8'hFF;
		16'hF840: out_word = 8'hFF;
		16'hF841: out_word = 8'hFF;
		16'hF842: out_word = 8'hFF;
		16'hF843: out_word = 8'hFF;
		16'hF844: out_word = 8'hFF;
		16'hF845: out_word = 8'hFF;
		16'hF846: out_word = 8'hFF;
		16'hF847: out_word = 8'hFF;
		16'hF848: out_word = 8'hFF;
		16'hF849: out_word = 8'hFF;
		16'hF84A: out_word = 8'hFF;
		16'hF84B: out_word = 8'hFF;
		16'hF84C: out_word = 8'hFF;
		16'hF84D: out_word = 8'hFF;
		16'hF84E: out_word = 8'hFF;
		16'hF84F: out_word = 8'hFF;
		16'hF850: out_word = 8'hFF;
		16'hF851: out_word = 8'hFF;
		16'hF852: out_word = 8'hFF;
		16'hF853: out_word = 8'hFF;
		16'hF854: out_word = 8'hFF;
		16'hF855: out_word = 8'hFF;
		16'hF856: out_word = 8'hFF;
		16'hF857: out_word = 8'hFF;
		16'hF858: out_word = 8'hFF;
		16'hF859: out_word = 8'hFF;
		16'hF85A: out_word = 8'hFF;
		16'hF85B: out_word = 8'hFF;
		16'hF85C: out_word = 8'hFF;
		16'hF85D: out_word = 8'hFF;
		16'hF85E: out_word = 8'hFF;
		16'hF85F: out_word = 8'hFF;
		16'hF860: out_word = 8'hFF;
		16'hF861: out_word = 8'hFF;
		16'hF862: out_word = 8'hFF;
		16'hF863: out_word = 8'hFF;
		16'hF864: out_word = 8'hFF;
		16'hF865: out_word = 8'hFF;
		16'hF866: out_word = 8'hFF;
		16'hF867: out_word = 8'hFF;
		16'hF868: out_word = 8'hFF;
		16'hF869: out_word = 8'hFF;
		16'hF86A: out_word = 8'hFF;
		16'hF86B: out_word = 8'hFF;
		16'hF86C: out_word = 8'hFF;
		16'hF86D: out_word = 8'hFF;
		16'hF86E: out_word = 8'hFF;
		16'hF86F: out_word = 8'hFF;
		16'hF870: out_word = 8'hFF;
		16'hF871: out_word = 8'hFF;
		16'hF872: out_word = 8'hFF;
		16'hF873: out_word = 8'hFF;
		16'hF874: out_word = 8'hFF;
		16'hF875: out_word = 8'hFF;
		16'hF876: out_word = 8'hFF;
		16'hF877: out_word = 8'hFF;
		16'hF878: out_word = 8'hFF;
		16'hF879: out_word = 8'hFF;
		16'hF87A: out_word = 8'hFF;
		16'hF87B: out_word = 8'hFF;
		16'hF87C: out_word = 8'hFF;
		16'hF87D: out_word = 8'hFF;
		16'hF87E: out_word = 8'hFF;
		16'hF87F: out_word = 8'hFF;
		16'hF880: out_word = 8'hFF;
		16'hF881: out_word = 8'hFF;
		16'hF882: out_word = 8'hFF;
		16'hF883: out_word = 8'hFF;
		16'hF884: out_word = 8'hFF;
		16'hF885: out_word = 8'hFF;
		16'hF886: out_word = 8'hFF;
		16'hF887: out_word = 8'hFF;
		16'hF888: out_word = 8'hFF;
		16'hF889: out_word = 8'hFF;
		16'hF88A: out_word = 8'hFF;
		16'hF88B: out_word = 8'hFF;
		16'hF88C: out_word = 8'hFF;
		16'hF88D: out_word = 8'hFF;
		16'hF88E: out_word = 8'hFF;
		16'hF88F: out_word = 8'hFF;
		16'hF890: out_word = 8'hFF;
		16'hF891: out_word = 8'hFF;
		16'hF892: out_word = 8'hFF;
		16'hF893: out_word = 8'hFF;
		16'hF894: out_word = 8'hFF;
		16'hF895: out_word = 8'hFF;
		16'hF896: out_word = 8'hFF;
		16'hF897: out_word = 8'hFF;
		16'hF898: out_word = 8'hFF;
		16'hF899: out_word = 8'hFF;
		16'hF89A: out_word = 8'hFF;
		16'hF89B: out_word = 8'hFF;
		16'hF89C: out_word = 8'hFF;
		16'hF89D: out_word = 8'hFF;
		16'hF89E: out_word = 8'hFF;
		16'hF89F: out_word = 8'hFF;
		16'hF8A0: out_word = 8'hFF;
		16'hF8A1: out_word = 8'hFF;
		16'hF8A2: out_word = 8'hFF;
		16'hF8A3: out_word = 8'hFF;
		16'hF8A4: out_word = 8'hFF;
		16'hF8A5: out_word = 8'hFF;
		16'hF8A6: out_word = 8'hFF;
		16'hF8A7: out_word = 8'hFF;
		16'hF8A8: out_word = 8'hFF;
		16'hF8A9: out_word = 8'hFF;
		16'hF8AA: out_word = 8'hFF;
		16'hF8AB: out_word = 8'hFF;
		16'hF8AC: out_word = 8'hFF;
		16'hF8AD: out_word = 8'hFF;
		16'hF8AE: out_word = 8'hFF;
		16'hF8AF: out_word = 8'hFF;
		16'hF8B0: out_word = 8'hFF;
		16'hF8B1: out_word = 8'hFF;
		16'hF8B2: out_word = 8'hFF;
		16'hF8B3: out_word = 8'hFF;
		16'hF8B4: out_word = 8'hFF;
		16'hF8B5: out_word = 8'hFF;
		16'hF8B6: out_word = 8'hFF;
		16'hF8B7: out_word = 8'hFF;
		16'hF8B8: out_word = 8'hFF;
		16'hF8B9: out_word = 8'hFF;
		16'hF8BA: out_word = 8'hFF;
		16'hF8BB: out_word = 8'hFF;
		16'hF8BC: out_word = 8'hFF;
		16'hF8BD: out_word = 8'hFF;
		16'hF8BE: out_word = 8'hFF;
		16'hF8BF: out_word = 8'hFF;
		16'hF8C0: out_word = 8'hFF;
		16'hF8C1: out_word = 8'hFF;
		16'hF8C2: out_word = 8'hFF;
		16'hF8C3: out_word = 8'hFF;
		16'hF8C4: out_word = 8'hFF;
		16'hF8C5: out_word = 8'hFF;
		16'hF8C6: out_word = 8'hFF;
		16'hF8C7: out_word = 8'hFF;
		16'hF8C8: out_word = 8'hFF;
		16'hF8C9: out_word = 8'hFF;
		16'hF8CA: out_word = 8'hFF;
		16'hF8CB: out_word = 8'hFF;
		16'hF8CC: out_word = 8'hFF;
		16'hF8CD: out_word = 8'hFF;
		16'hF8CE: out_word = 8'hFF;
		16'hF8CF: out_word = 8'hFF;
		16'hF8D0: out_word = 8'hFF;
		16'hF8D1: out_word = 8'hFF;
		16'hF8D2: out_word = 8'hFF;
		16'hF8D3: out_word = 8'hFF;
		16'hF8D4: out_word = 8'hFF;
		16'hF8D5: out_word = 8'hFF;
		16'hF8D6: out_word = 8'hFF;
		16'hF8D7: out_word = 8'hFF;
		16'hF8D8: out_word = 8'hFF;
		16'hF8D9: out_word = 8'hFF;
		16'hF8DA: out_word = 8'hFF;
		16'hF8DB: out_word = 8'hFF;
		16'hF8DC: out_word = 8'hFF;
		16'hF8DD: out_word = 8'hFF;
		16'hF8DE: out_word = 8'hFF;
		16'hF8DF: out_word = 8'hFF;
		16'hF8E0: out_word = 8'hFF;
		16'hF8E1: out_word = 8'hFF;
		16'hF8E2: out_word = 8'hFF;
		16'hF8E3: out_word = 8'hFF;
		16'hF8E4: out_word = 8'hFF;
		16'hF8E5: out_word = 8'hFF;
		16'hF8E6: out_word = 8'hFF;
		16'hF8E7: out_word = 8'hFF;
		16'hF8E8: out_word = 8'hFF;
		16'hF8E9: out_word = 8'hFF;
		16'hF8EA: out_word = 8'hFF;
		16'hF8EB: out_word = 8'hFF;
		16'hF8EC: out_word = 8'hFF;
		16'hF8ED: out_word = 8'hFF;
		16'hF8EE: out_word = 8'hFF;
		16'hF8EF: out_word = 8'hFF;
		16'hF8F0: out_word = 8'hFF;
		16'hF8F1: out_word = 8'hFF;
		16'hF8F2: out_word = 8'hFF;
		16'hF8F3: out_word = 8'hFF;
		16'hF8F4: out_word = 8'hFF;
		16'hF8F5: out_word = 8'hFF;
		16'hF8F6: out_word = 8'hFF;
		16'hF8F7: out_word = 8'hFF;
		16'hF8F8: out_word = 8'hFF;
		16'hF8F9: out_word = 8'hFF;
		16'hF8FA: out_word = 8'hFF;
		16'hF8FB: out_word = 8'hFF;
		16'hF8FC: out_word = 8'hFF;
		16'hF8FD: out_word = 8'hFF;
		16'hF8FE: out_word = 8'hFF;
		16'hF8FF: out_word = 8'hFF;
		16'hF900: out_word = 8'hFF;
		16'hF901: out_word = 8'hFF;
		16'hF902: out_word = 8'hFF;
		16'hF903: out_word = 8'hFF;
		16'hF904: out_word = 8'hFF;
		16'hF905: out_word = 8'hFF;
		16'hF906: out_word = 8'hFF;
		16'hF907: out_word = 8'hFF;
		16'hF908: out_word = 8'hFF;
		16'hF909: out_word = 8'hFF;
		16'hF90A: out_word = 8'hFF;
		16'hF90B: out_word = 8'hFF;
		16'hF90C: out_word = 8'hFF;
		16'hF90D: out_word = 8'hFF;
		16'hF90E: out_word = 8'hFF;
		16'hF90F: out_word = 8'hFF;
		16'hF910: out_word = 8'hFF;
		16'hF911: out_word = 8'hFF;
		16'hF912: out_word = 8'hFF;
		16'hF913: out_word = 8'hFF;
		16'hF914: out_word = 8'hFF;
		16'hF915: out_word = 8'hFF;
		16'hF916: out_word = 8'hFF;
		16'hF917: out_word = 8'hFF;
		16'hF918: out_word = 8'hFF;
		16'hF919: out_word = 8'hFF;
		16'hF91A: out_word = 8'hFF;
		16'hF91B: out_word = 8'hFF;
		16'hF91C: out_word = 8'hFF;
		16'hF91D: out_word = 8'hFF;
		16'hF91E: out_word = 8'hFF;
		16'hF91F: out_word = 8'hFF;
		16'hF920: out_word = 8'hFF;
		16'hF921: out_word = 8'hFF;
		16'hF922: out_word = 8'hFF;
		16'hF923: out_word = 8'hFF;
		16'hF924: out_word = 8'hFF;
		16'hF925: out_word = 8'hFF;
		16'hF926: out_word = 8'hFF;
		16'hF927: out_word = 8'hFF;
		16'hF928: out_word = 8'hFF;
		16'hF929: out_word = 8'hFF;
		16'hF92A: out_word = 8'hFF;
		16'hF92B: out_word = 8'hFF;
		16'hF92C: out_word = 8'hFF;
		16'hF92D: out_word = 8'hFF;
		16'hF92E: out_word = 8'hFF;
		16'hF92F: out_word = 8'hFF;
		16'hF930: out_word = 8'hFF;
		16'hF931: out_word = 8'hFF;
		16'hF932: out_word = 8'hFF;
		16'hF933: out_word = 8'hFF;
		16'hF934: out_word = 8'hFF;
		16'hF935: out_word = 8'hFF;
		16'hF936: out_word = 8'hFF;
		16'hF937: out_word = 8'hFF;
		16'hF938: out_word = 8'hFF;
		16'hF939: out_word = 8'hFF;
		16'hF93A: out_word = 8'hFF;
		16'hF93B: out_word = 8'hFF;
		16'hF93C: out_word = 8'hFF;
		16'hF93D: out_word = 8'hFF;
		16'hF93E: out_word = 8'hFF;
		16'hF93F: out_word = 8'hFF;
		16'hF940: out_word = 8'hFF;
		16'hF941: out_word = 8'hFF;
		16'hF942: out_word = 8'hFF;
		16'hF943: out_word = 8'hFF;
		16'hF944: out_word = 8'hFF;
		16'hF945: out_word = 8'hFF;
		16'hF946: out_word = 8'hFF;
		16'hF947: out_word = 8'hFF;
		16'hF948: out_word = 8'hFF;
		16'hF949: out_word = 8'hFF;
		16'hF94A: out_word = 8'hFF;
		16'hF94B: out_word = 8'hFF;
		16'hF94C: out_word = 8'hFF;
		16'hF94D: out_word = 8'hFF;
		16'hF94E: out_word = 8'hFF;
		16'hF94F: out_word = 8'hFF;
		16'hF950: out_word = 8'hFF;
		16'hF951: out_word = 8'hFF;
		16'hF952: out_word = 8'hFF;
		16'hF953: out_word = 8'hFF;
		16'hF954: out_word = 8'hFF;
		16'hF955: out_word = 8'hFF;
		16'hF956: out_word = 8'hFF;
		16'hF957: out_word = 8'hFF;
		16'hF958: out_word = 8'hFF;
		16'hF959: out_word = 8'hFF;
		16'hF95A: out_word = 8'hFF;
		16'hF95B: out_word = 8'hFF;
		16'hF95C: out_word = 8'hFF;
		16'hF95D: out_word = 8'hFF;
		16'hF95E: out_word = 8'hFF;
		16'hF95F: out_word = 8'hFF;
		16'hF960: out_word = 8'hFF;
		16'hF961: out_word = 8'hFF;
		16'hF962: out_word = 8'hFF;
		16'hF963: out_word = 8'hFF;
		16'hF964: out_word = 8'hFF;
		16'hF965: out_word = 8'hFF;
		16'hF966: out_word = 8'hFF;
		16'hF967: out_word = 8'hFF;
		16'hF968: out_word = 8'hFF;
		16'hF969: out_word = 8'hFF;
		16'hF96A: out_word = 8'hFF;
		16'hF96B: out_word = 8'hFF;
		16'hF96C: out_word = 8'hFF;
		16'hF96D: out_word = 8'hFF;
		16'hF96E: out_word = 8'hFF;
		16'hF96F: out_word = 8'hFF;
		16'hF970: out_word = 8'hFF;
		16'hF971: out_word = 8'hFF;
		16'hF972: out_word = 8'hFF;
		16'hF973: out_word = 8'hFF;
		16'hF974: out_word = 8'hFF;
		16'hF975: out_word = 8'hFF;
		16'hF976: out_word = 8'hFF;
		16'hF977: out_word = 8'hFF;
		16'hF978: out_word = 8'hFF;
		16'hF979: out_word = 8'hFF;
		16'hF97A: out_word = 8'hFF;
		16'hF97B: out_word = 8'hFF;
		16'hF97C: out_word = 8'hFF;
		16'hF97D: out_word = 8'hFF;
		16'hF97E: out_word = 8'hFF;
		16'hF97F: out_word = 8'hFF;
		16'hF980: out_word = 8'hFF;
		16'hF981: out_word = 8'hFF;
		16'hF982: out_word = 8'hFF;
		16'hF983: out_word = 8'hFF;
		16'hF984: out_word = 8'hFF;
		16'hF985: out_word = 8'hFF;
		16'hF986: out_word = 8'hFF;
		16'hF987: out_word = 8'hFF;
		16'hF988: out_word = 8'hFF;
		16'hF989: out_word = 8'hFF;
		16'hF98A: out_word = 8'hFF;
		16'hF98B: out_word = 8'hFF;
		16'hF98C: out_word = 8'hFF;
		16'hF98D: out_word = 8'hFF;
		16'hF98E: out_word = 8'hFF;
		16'hF98F: out_word = 8'hFF;
		16'hF990: out_word = 8'hFF;
		16'hF991: out_word = 8'hFF;
		16'hF992: out_word = 8'hFF;
		16'hF993: out_word = 8'hFF;
		16'hF994: out_word = 8'hFF;
		16'hF995: out_word = 8'hFF;
		16'hF996: out_word = 8'hFF;
		16'hF997: out_word = 8'hFF;
		16'hF998: out_word = 8'hFF;
		16'hF999: out_word = 8'hFF;
		16'hF99A: out_word = 8'hFF;
		16'hF99B: out_word = 8'hFF;
		16'hF99C: out_word = 8'hFF;
		16'hF99D: out_word = 8'hFF;
		16'hF99E: out_word = 8'hFF;
		16'hF99F: out_word = 8'hFF;
		16'hF9A0: out_word = 8'hFF;
		16'hF9A1: out_word = 8'hFF;
		16'hF9A2: out_word = 8'hFF;
		16'hF9A3: out_word = 8'hFF;
		16'hF9A4: out_word = 8'hFF;
		16'hF9A5: out_word = 8'hFF;
		16'hF9A6: out_word = 8'hFF;
		16'hF9A7: out_word = 8'hFF;
		16'hF9A8: out_word = 8'hFF;
		16'hF9A9: out_word = 8'hFF;
		16'hF9AA: out_word = 8'hFF;
		16'hF9AB: out_word = 8'hFF;
		16'hF9AC: out_word = 8'hFF;
		16'hF9AD: out_word = 8'hFF;
		16'hF9AE: out_word = 8'hFF;
		16'hF9AF: out_word = 8'hFF;
		16'hF9B0: out_word = 8'hFF;
		16'hF9B1: out_word = 8'hFF;
		16'hF9B2: out_word = 8'hFF;
		16'hF9B3: out_word = 8'hFF;
		16'hF9B4: out_word = 8'hFF;
		16'hF9B5: out_word = 8'hFF;
		16'hF9B6: out_word = 8'hFF;
		16'hF9B7: out_word = 8'hFF;
		16'hF9B8: out_word = 8'hFF;
		16'hF9B9: out_word = 8'hFF;
		16'hF9BA: out_word = 8'hFF;
		16'hF9BB: out_word = 8'hFF;
		16'hF9BC: out_word = 8'hFF;
		16'hF9BD: out_word = 8'hFF;
		16'hF9BE: out_word = 8'hFF;
		16'hF9BF: out_word = 8'hFF;
		16'hF9C0: out_word = 8'hFF;
		16'hF9C1: out_word = 8'hFF;
		16'hF9C2: out_word = 8'hFF;
		16'hF9C3: out_word = 8'hFF;
		16'hF9C4: out_word = 8'hFF;
		16'hF9C5: out_word = 8'hFF;
		16'hF9C6: out_word = 8'hFF;
		16'hF9C7: out_word = 8'hFF;
		16'hF9C8: out_word = 8'hFF;
		16'hF9C9: out_word = 8'hFF;
		16'hF9CA: out_word = 8'hFF;
		16'hF9CB: out_word = 8'hFF;
		16'hF9CC: out_word = 8'hFF;
		16'hF9CD: out_word = 8'hFF;
		16'hF9CE: out_word = 8'hFF;
		16'hF9CF: out_word = 8'hFF;
		16'hF9D0: out_word = 8'hFF;
		16'hF9D1: out_word = 8'hFF;
		16'hF9D2: out_word = 8'hFF;
		16'hF9D3: out_word = 8'hFF;
		16'hF9D4: out_word = 8'hFF;
		16'hF9D5: out_word = 8'hFF;
		16'hF9D6: out_word = 8'hFF;
		16'hF9D7: out_word = 8'hFF;
		16'hF9D8: out_word = 8'hFF;
		16'hF9D9: out_word = 8'hFF;
		16'hF9DA: out_word = 8'hFF;
		16'hF9DB: out_word = 8'hFF;
		16'hF9DC: out_word = 8'hFF;
		16'hF9DD: out_word = 8'hFF;
		16'hF9DE: out_word = 8'hFF;
		16'hF9DF: out_word = 8'hFF;
		16'hF9E0: out_word = 8'hFF;
		16'hF9E1: out_word = 8'hFF;
		16'hF9E2: out_word = 8'hFF;
		16'hF9E3: out_word = 8'hFF;
		16'hF9E4: out_word = 8'hFF;
		16'hF9E5: out_word = 8'hFF;
		16'hF9E6: out_word = 8'hFF;
		16'hF9E7: out_word = 8'hFF;
		16'hF9E8: out_word = 8'hFF;
		16'hF9E9: out_word = 8'hFF;
		16'hF9EA: out_word = 8'hFF;
		16'hF9EB: out_word = 8'hFF;
		16'hF9EC: out_word = 8'hFF;
		16'hF9ED: out_word = 8'hFF;
		16'hF9EE: out_word = 8'hFF;
		16'hF9EF: out_word = 8'hFF;
		16'hF9F0: out_word = 8'hFF;
		16'hF9F1: out_word = 8'hFF;
		16'hF9F2: out_word = 8'hFF;
		16'hF9F3: out_word = 8'hFF;
		16'hF9F4: out_word = 8'hFF;
		16'hF9F5: out_word = 8'hFF;
		16'hF9F6: out_word = 8'hFF;
		16'hF9F7: out_word = 8'hFF;
		16'hF9F8: out_word = 8'hFF;
		16'hF9F9: out_word = 8'hFF;
		16'hF9FA: out_word = 8'hFF;
		16'hF9FB: out_word = 8'hFF;
		16'hF9FC: out_word = 8'hFF;
		16'hF9FD: out_word = 8'hFF;
		16'hF9FE: out_word = 8'hFF;
		16'hF9FF: out_word = 8'hFF;
		16'hFA00: out_word = 8'hFF;
		16'hFA01: out_word = 8'hFF;
		16'hFA02: out_word = 8'hFF;
		16'hFA03: out_word = 8'hFF;
		16'hFA04: out_word = 8'hFF;
		16'hFA05: out_word = 8'hFF;
		16'hFA06: out_word = 8'hFF;
		16'hFA07: out_word = 8'hFF;
		16'hFA08: out_word = 8'hFF;
		16'hFA09: out_word = 8'hFF;
		16'hFA0A: out_word = 8'hFF;
		16'hFA0B: out_word = 8'hFF;
		16'hFA0C: out_word = 8'hFF;
		16'hFA0D: out_word = 8'hFF;
		16'hFA0E: out_word = 8'hFF;
		16'hFA0F: out_word = 8'hFF;
		16'hFA10: out_word = 8'hFF;
		16'hFA11: out_word = 8'hFF;
		16'hFA12: out_word = 8'hFF;
		16'hFA13: out_word = 8'hFF;
		16'hFA14: out_word = 8'hFF;
		16'hFA15: out_word = 8'hFF;
		16'hFA16: out_word = 8'hFF;
		16'hFA17: out_word = 8'hFF;
		16'hFA18: out_word = 8'hFF;
		16'hFA19: out_word = 8'hFF;
		16'hFA1A: out_word = 8'hFF;
		16'hFA1B: out_word = 8'hFF;
		16'hFA1C: out_word = 8'hFF;
		16'hFA1D: out_word = 8'hFF;
		16'hFA1E: out_word = 8'hFF;
		16'hFA1F: out_word = 8'hFF;
		16'hFA20: out_word = 8'hFF;
		16'hFA21: out_word = 8'hFF;
		16'hFA22: out_word = 8'hFF;
		16'hFA23: out_word = 8'hFF;
		16'hFA24: out_word = 8'hFF;
		16'hFA25: out_word = 8'hFF;
		16'hFA26: out_word = 8'hFF;
		16'hFA27: out_word = 8'hFF;
		16'hFA28: out_word = 8'hFF;
		16'hFA29: out_word = 8'hFF;
		16'hFA2A: out_word = 8'hFF;
		16'hFA2B: out_word = 8'hFF;
		16'hFA2C: out_word = 8'hFF;
		16'hFA2D: out_word = 8'hFF;
		16'hFA2E: out_word = 8'hFF;
		16'hFA2F: out_word = 8'hFF;
		16'hFA30: out_word = 8'hFF;
		16'hFA31: out_word = 8'hFF;
		16'hFA32: out_word = 8'hFF;
		16'hFA33: out_word = 8'hFF;
		16'hFA34: out_word = 8'hFF;
		16'hFA35: out_word = 8'hFF;
		16'hFA36: out_word = 8'hFF;
		16'hFA37: out_word = 8'hFF;
		16'hFA38: out_word = 8'hFF;
		16'hFA39: out_word = 8'hFF;
		16'hFA3A: out_word = 8'hFF;
		16'hFA3B: out_word = 8'hFF;
		16'hFA3C: out_word = 8'hFF;
		16'hFA3D: out_word = 8'hFF;
		16'hFA3E: out_word = 8'hFF;
		16'hFA3F: out_word = 8'hFF;
		16'hFA40: out_word = 8'hFF;
		16'hFA41: out_word = 8'hFF;
		16'hFA42: out_word = 8'hFF;
		16'hFA43: out_word = 8'hFF;
		16'hFA44: out_word = 8'hFF;
		16'hFA45: out_word = 8'hFF;
		16'hFA46: out_word = 8'hFF;
		16'hFA47: out_word = 8'hFF;
		16'hFA48: out_word = 8'hFF;
		16'hFA49: out_word = 8'hFF;
		16'hFA4A: out_word = 8'hFF;
		16'hFA4B: out_word = 8'hFF;
		16'hFA4C: out_word = 8'hFF;
		16'hFA4D: out_word = 8'hFF;
		16'hFA4E: out_word = 8'hFF;
		16'hFA4F: out_word = 8'hFF;
		16'hFA50: out_word = 8'hFF;
		16'hFA51: out_word = 8'hFF;
		16'hFA52: out_word = 8'hFF;
		16'hFA53: out_word = 8'hFF;
		16'hFA54: out_word = 8'hFF;
		16'hFA55: out_word = 8'hFF;
		16'hFA56: out_word = 8'hFF;
		16'hFA57: out_word = 8'hFF;
		16'hFA58: out_word = 8'hFF;
		16'hFA59: out_word = 8'hFF;
		16'hFA5A: out_word = 8'hFF;
		16'hFA5B: out_word = 8'hFF;
		16'hFA5C: out_word = 8'hFF;
		16'hFA5D: out_word = 8'hFF;
		16'hFA5E: out_word = 8'hFF;
		16'hFA5F: out_word = 8'hFF;
		16'hFA60: out_word = 8'hFF;
		16'hFA61: out_word = 8'hFF;
		16'hFA62: out_word = 8'hFF;
		16'hFA63: out_word = 8'hFF;
		16'hFA64: out_word = 8'hFF;
		16'hFA65: out_word = 8'hFF;
		16'hFA66: out_word = 8'hFF;
		16'hFA67: out_word = 8'hFF;
		16'hFA68: out_word = 8'hFF;
		16'hFA69: out_word = 8'hFF;
		16'hFA6A: out_word = 8'hFF;
		16'hFA6B: out_word = 8'hFF;
		16'hFA6C: out_word = 8'hFF;
		16'hFA6D: out_word = 8'hFF;
		16'hFA6E: out_word = 8'hFF;
		16'hFA6F: out_word = 8'hFF;
		16'hFA70: out_word = 8'hFF;
		16'hFA71: out_word = 8'hFF;
		16'hFA72: out_word = 8'hFF;
		16'hFA73: out_word = 8'hFF;
		16'hFA74: out_word = 8'hFF;
		16'hFA75: out_word = 8'hFF;
		16'hFA76: out_word = 8'hFF;
		16'hFA77: out_word = 8'hFF;
		16'hFA78: out_word = 8'hFF;
		16'hFA79: out_word = 8'hFF;
		16'hFA7A: out_word = 8'hFF;
		16'hFA7B: out_word = 8'hFF;
		16'hFA7C: out_word = 8'hFF;
		16'hFA7D: out_word = 8'hFF;
		16'hFA7E: out_word = 8'hFF;
		16'hFA7F: out_word = 8'hFF;
		16'hFA80: out_word = 8'hFF;
		16'hFA81: out_word = 8'hFF;
		16'hFA82: out_word = 8'hFF;
		16'hFA83: out_word = 8'hFF;
		16'hFA84: out_word = 8'hFF;
		16'hFA85: out_word = 8'hFF;
		16'hFA86: out_word = 8'hFF;
		16'hFA87: out_word = 8'hFF;
		16'hFA88: out_word = 8'hFF;
		16'hFA89: out_word = 8'hFF;
		16'hFA8A: out_word = 8'hFF;
		16'hFA8B: out_word = 8'hFF;
		16'hFA8C: out_word = 8'hFF;
		16'hFA8D: out_word = 8'hFF;
		16'hFA8E: out_word = 8'hFF;
		16'hFA8F: out_word = 8'hFF;
		16'hFA90: out_word = 8'hFF;
		16'hFA91: out_word = 8'hFF;
		16'hFA92: out_word = 8'hFF;
		16'hFA93: out_word = 8'hFF;
		16'hFA94: out_word = 8'hFF;
		16'hFA95: out_word = 8'hFF;
		16'hFA96: out_word = 8'hFF;
		16'hFA97: out_word = 8'hFF;
		16'hFA98: out_word = 8'hFF;
		16'hFA99: out_word = 8'hFF;
		16'hFA9A: out_word = 8'hFF;
		16'hFA9B: out_word = 8'hFF;
		16'hFA9C: out_word = 8'hFF;
		16'hFA9D: out_word = 8'hFF;
		16'hFA9E: out_word = 8'hFF;
		16'hFA9F: out_word = 8'hFF;
		16'hFAA0: out_word = 8'hFF;
		16'hFAA1: out_word = 8'hFF;
		16'hFAA2: out_word = 8'hFF;
		16'hFAA3: out_word = 8'hFF;
		16'hFAA4: out_word = 8'hFF;
		16'hFAA5: out_word = 8'hFF;
		16'hFAA6: out_word = 8'hFF;
		16'hFAA7: out_word = 8'hFF;
		16'hFAA8: out_word = 8'hFF;
		16'hFAA9: out_word = 8'hFF;
		16'hFAAA: out_word = 8'hFF;
		16'hFAAB: out_word = 8'hFF;
		16'hFAAC: out_word = 8'hFF;
		16'hFAAD: out_word = 8'hFF;
		16'hFAAE: out_word = 8'hFF;
		16'hFAAF: out_word = 8'hFF;
		16'hFAB0: out_word = 8'hFF;
		16'hFAB1: out_word = 8'hFF;
		16'hFAB2: out_word = 8'hFF;
		16'hFAB3: out_word = 8'hFF;
		16'hFAB4: out_word = 8'hFF;
		16'hFAB5: out_word = 8'hFF;
		16'hFAB6: out_word = 8'hFF;
		16'hFAB7: out_word = 8'hFF;
		16'hFAB8: out_word = 8'hFF;
		16'hFAB9: out_word = 8'hFF;
		16'hFABA: out_word = 8'hFF;
		16'hFABB: out_word = 8'hFF;
		16'hFABC: out_word = 8'hFF;
		16'hFABD: out_word = 8'hFF;
		16'hFABE: out_word = 8'hFF;
		16'hFABF: out_word = 8'hFF;
		16'hFAC0: out_word = 8'hFF;
		16'hFAC1: out_word = 8'hFF;
		16'hFAC2: out_word = 8'hFF;
		16'hFAC3: out_word = 8'hFF;
		16'hFAC4: out_word = 8'hFF;
		16'hFAC5: out_word = 8'hFF;
		16'hFAC6: out_word = 8'hFF;
		16'hFAC7: out_word = 8'hFF;
		16'hFAC8: out_word = 8'hFF;
		16'hFAC9: out_word = 8'hFF;
		16'hFACA: out_word = 8'hFF;
		16'hFACB: out_word = 8'hFF;
		16'hFACC: out_word = 8'hFF;
		16'hFACD: out_word = 8'hFF;
		16'hFACE: out_word = 8'hFF;
		16'hFACF: out_word = 8'hFF;
		16'hFAD0: out_word = 8'hFF;
		16'hFAD1: out_word = 8'hFF;
		16'hFAD2: out_word = 8'hFF;
		16'hFAD3: out_word = 8'hFF;
		16'hFAD4: out_word = 8'hFF;
		16'hFAD5: out_word = 8'hFF;
		16'hFAD6: out_word = 8'hFF;
		16'hFAD7: out_word = 8'hFF;
		16'hFAD8: out_word = 8'hFF;
		16'hFAD9: out_word = 8'hFF;
		16'hFADA: out_word = 8'hFF;
		16'hFADB: out_word = 8'hFF;
		16'hFADC: out_word = 8'hFF;
		16'hFADD: out_word = 8'hFF;
		16'hFADE: out_word = 8'hFF;
		16'hFADF: out_word = 8'hFF;
		16'hFAE0: out_word = 8'hFF;
		16'hFAE1: out_word = 8'hFF;
		16'hFAE2: out_word = 8'hFF;
		16'hFAE3: out_word = 8'hFF;
		16'hFAE4: out_word = 8'hFF;
		16'hFAE5: out_word = 8'hFF;
		16'hFAE6: out_word = 8'hFF;
		16'hFAE7: out_word = 8'hFF;
		16'hFAE8: out_word = 8'hFF;
		16'hFAE9: out_word = 8'hFF;
		16'hFAEA: out_word = 8'hFF;
		16'hFAEB: out_word = 8'hFF;
		16'hFAEC: out_word = 8'hFF;
		16'hFAED: out_word = 8'hFF;
		16'hFAEE: out_word = 8'hFF;
		16'hFAEF: out_word = 8'hFF;
		16'hFAF0: out_word = 8'hFF;
		16'hFAF1: out_word = 8'hFF;
		16'hFAF2: out_word = 8'hFF;
		16'hFAF3: out_word = 8'hFF;
		16'hFAF4: out_word = 8'hFF;
		16'hFAF5: out_word = 8'hFF;
		16'hFAF6: out_word = 8'hFF;
		16'hFAF7: out_word = 8'hFF;
		16'hFAF8: out_word = 8'hFF;
		16'hFAF9: out_word = 8'hFF;
		16'hFAFA: out_word = 8'hFF;
		16'hFAFB: out_word = 8'hFF;
		16'hFAFC: out_word = 8'hFF;
		16'hFAFD: out_word = 8'hFF;
		16'hFAFE: out_word = 8'hFF;
		16'hFAFF: out_word = 8'hFF;
		16'hFB00: out_word = 8'hFF;
		16'hFB01: out_word = 8'hFF;
		16'hFB02: out_word = 8'hFF;
		16'hFB03: out_word = 8'hFF;
		16'hFB04: out_word = 8'hFF;
		16'hFB05: out_word = 8'hFF;
		16'hFB06: out_word = 8'hFF;
		16'hFB07: out_word = 8'hFF;
		16'hFB08: out_word = 8'hFF;
		16'hFB09: out_word = 8'hFF;
		16'hFB0A: out_word = 8'hFF;
		16'hFB0B: out_word = 8'hFF;
		16'hFB0C: out_word = 8'hFF;
		16'hFB0D: out_word = 8'hFF;
		16'hFB0E: out_word = 8'hFF;
		16'hFB0F: out_word = 8'hFF;
		16'hFB10: out_word = 8'hFF;
		16'hFB11: out_word = 8'hFF;
		16'hFB12: out_word = 8'hFF;
		16'hFB13: out_word = 8'hFF;
		16'hFB14: out_word = 8'hFF;
		16'hFB15: out_word = 8'hFF;
		16'hFB16: out_word = 8'hFF;
		16'hFB17: out_word = 8'hFF;
		16'hFB18: out_word = 8'hFF;
		16'hFB19: out_word = 8'hFF;
		16'hFB1A: out_word = 8'hFF;
		16'hFB1B: out_word = 8'hFF;
		16'hFB1C: out_word = 8'hFF;
		16'hFB1D: out_word = 8'hFF;
		16'hFB1E: out_word = 8'hFF;
		16'hFB1F: out_word = 8'hFF;
		16'hFB20: out_word = 8'hFF;
		16'hFB21: out_word = 8'hFF;
		16'hFB22: out_word = 8'hFF;
		16'hFB23: out_word = 8'hFF;
		16'hFB24: out_word = 8'hFF;
		16'hFB25: out_word = 8'hFF;
		16'hFB26: out_word = 8'hFF;
		16'hFB27: out_word = 8'hFF;
		16'hFB28: out_word = 8'hFF;
		16'hFB29: out_word = 8'hFF;
		16'hFB2A: out_word = 8'hFF;
		16'hFB2B: out_word = 8'hFF;
		16'hFB2C: out_word = 8'hFF;
		16'hFB2D: out_word = 8'hFF;
		16'hFB2E: out_word = 8'hFF;
		16'hFB2F: out_word = 8'hFF;
		16'hFB30: out_word = 8'hFF;
		16'hFB31: out_word = 8'hFF;
		16'hFB32: out_word = 8'hFF;
		16'hFB33: out_word = 8'hFF;
		16'hFB34: out_word = 8'hFF;
		16'hFB35: out_word = 8'hFF;
		16'hFB36: out_word = 8'hFF;
		16'hFB37: out_word = 8'hFF;
		16'hFB38: out_word = 8'hFF;
		16'hFB39: out_word = 8'hFF;
		16'hFB3A: out_word = 8'hFF;
		16'hFB3B: out_word = 8'hFF;
		16'hFB3C: out_word = 8'hFF;
		16'hFB3D: out_word = 8'hFF;
		16'hFB3E: out_word = 8'hFF;
		16'hFB3F: out_word = 8'hFF;
		16'hFB40: out_word = 8'hFF;
		16'hFB41: out_word = 8'hFF;
		16'hFB42: out_word = 8'hFF;
		16'hFB43: out_word = 8'hFF;
		16'hFB44: out_word = 8'hFF;
		16'hFB45: out_word = 8'hFF;
		16'hFB46: out_word = 8'hFF;
		16'hFB47: out_word = 8'hFF;
		16'hFB48: out_word = 8'hFF;
		16'hFB49: out_word = 8'hFF;
		16'hFB4A: out_word = 8'hFF;
		16'hFB4B: out_word = 8'hFF;
		16'hFB4C: out_word = 8'hFF;
		16'hFB4D: out_word = 8'hFF;
		16'hFB4E: out_word = 8'hFF;
		16'hFB4F: out_word = 8'hFF;
		16'hFB50: out_word = 8'hFF;
		16'hFB51: out_word = 8'hFF;
		16'hFB52: out_word = 8'hFF;
		16'hFB53: out_word = 8'hFF;
		16'hFB54: out_word = 8'hFF;
		16'hFB55: out_word = 8'hFF;
		16'hFB56: out_word = 8'hFF;
		16'hFB57: out_word = 8'hFF;
		16'hFB58: out_word = 8'hFF;
		16'hFB59: out_word = 8'hFF;
		16'hFB5A: out_word = 8'hFF;
		16'hFB5B: out_word = 8'hFF;
		16'hFB5C: out_word = 8'hFF;
		16'hFB5D: out_word = 8'hFF;
		16'hFB5E: out_word = 8'hFF;
		16'hFB5F: out_word = 8'hFF;
		16'hFB60: out_word = 8'hFF;
		16'hFB61: out_word = 8'hFF;
		16'hFB62: out_word = 8'hFF;
		16'hFB63: out_word = 8'hFF;
		16'hFB64: out_word = 8'hFF;
		16'hFB65: out_word = 8'hFF;
		16'hFB66: out_word = 8'hFF;
		16'hFB67: out_word = 8'hFF;
		16'hFB68: out_word = 8'hFF;
		16'hFB69: out_word = 8'hFF;
		16'hFB6A: out_word = 8'hFF;
		16'hFB6B: out_word = 8'hFF;
		16'hFB6C: out_word = 8'hFF;
		16'hFB6D: out_word = 8'hFF;
		16'hFB6E: out_word = 8'hFF;
		16'hFB6F: out_word = 8'hFF;
		16'hFB70: out_word = 8'hFF;
		16'hFB71: out_word = 8'hFF;
		16'hFB72: out_word = 8'hFF;
		16'hFB73: out_word = 8'hFF;
		16'hFB74: out_word = 8'hFF;
		16'hFB75: out_word = 8'hFF;
		16'hFB76: out_word = 8'hFF;
		16'hFB77: out_word = 8'hFF;
		16'hFB78: out_word = 8'hFF;
		16'hFB79: out_word = 8'hFF;
		16'hFB7A: out_word = 8'hFF;
		16'hFB7B: out_word = 8'hFF;
		16'hFB7C: out_word = 8'hFF;
		16'hFB7D: out_word = 8'hFF;
		16'hFB7E: out_word = 8'hFF;
		16'hFB7F: out_word = 8'hFF;
		16'hFB80: out_word = 8'hFF;
		16'hFB81: out_word = 8'hFF;
		16'hFB82: out_word = 8'hFF;
		16'hFB83: out_word = 8'hFF;
		16'hFB84: out_word = 8'hFF;
		16'hFB85: out_word = 8'hFF;
		16'hFB86: out_word = 8'hFF;
		16'hFB87: out_word = 8'hFF;
		16'hFB88: out_word = 8'hFF;
		16'hFB89: out_word = 8'hFF;
		16'hFB8A: out_word = 8'hFF;
		16'hFB8B: out_word = 8'hFF;
		16'hFB8C: out_word = 8'hFF;
		16'hFB8D: out_word = 8'hFF;
		16'hFB8E: out_word = 8'hFF;
		16'hFB8F: out_word = 8'hFF;
		16'hFB90: out_word = 8'hFF;
		16'hFB91: out_word = 8'hFF;
		16'hFB92: out_word = 8'hFF;
		16'hFB93: out_word = 8'hFF;
		16'hFB94: out_word = 8'hFF;
		16'hFB95: out_word = 8'hFF;
		16'hFB96: out_word = 8'hFF;
		16'hFB97: out_word = 8'hFF;
		16'hFB98: out_word = 8'hFF;
		16'hFB99: out_word = 8'hFF;
		16'hFB9A: out_word = 8'hFF;
		16'hFB9B: out_word = 8'hFF;
		16'hFB9C: out_word = 8'hFF;
		16'hFB9D: out_word = 8'hFF;
		16'hFB9E: out_word = 8'hFF;
		16'hFB9F: out_word = 8'hFF;
		16'hFBA0: out_word = 8'hFF;
		16'hFBA1: out_word = 8'hFF;
		16'hFBA2: out_word = 8'hFF;
		16'hFBA3: out_word = 8'hFF;
		16'hFBA4: out_word = 8'hFF;
		16'hFBA5: out_word = 8'hFF;
		16'hFBA6: out_word = 8'hFF;
		16'hFBA7: out_word = 8'hFF;
		16'hFBA8: out_word = 8'hFF;
		16'hFBA9: out_word = 8'hFF;
		16'hFBAA: out_word = 8'hFF;
		16'hFBAB: out_word = 8'hFF;
		16'hFBAC: out_word = 8'hFF;
		16'hFBAD: out_word = 8'hFF;
		16'hFBAE: out_word = 8'hFF;
		16'hFBAF: out_word = 8'hFF;
		16'hFBB0: out_word = 8'hFF;
		16'hFBB1: out_word = 8'hFF;
		16'hFBB2: out_word = 8'hFF;
		16'hFBB3: out_word = 8'hFF;
		16'hFBB4: out_word = 8'hFF;
		16'hFBB5: out_word = 8'hFF;
		16'hFBB6: out_word = 8'hFF;
		16'hFBB7: out_word = 8'hFF;
		16'hFBB8: out_word = 8'hFF;
		16'hFBB9: out_word = 8'hFF;
		16'hFBBA: out_word = 8'hFF;
		16'hFBBB: out_word = 8'hFF;
		16'hFBBC: out_word = 8'hFF;
		16'hFBBD: out_word = 8'hFF;
		16'hFBBE: out_word = 8'hFF;
		16'hFBBF: out_word = 8'hFF;
		16'hFBC0: out_word = 8'hFF;
		16'hFBC1: out_word = 8'hFF;
		16'hFBC2: out_word = 8'hFF;
		16'hFBC3: out_word = 8'hFF;
		16'hFBC4: out_word = 8'hFF;
		16'hFBC5: out_word = 8'hFF;
		16'hFBC6: out_word = 8'hFF;
		16'hFBC7: out_word = 8'hFF;
		16'hFBC8: out_word = 8'hFF;
		16'hFBC9: out_word = 8'hFF;
		16'hFBCA: out_word = 8'hFF;
		16'hFBCB: out_word = 8'hFF;
		16'hFBCC: out_word = 8'hFF;
		16'hFBCD: out_word = 8'hFF;
		16'hFBCE: out_word = 8'hFF;
		16'hFBCF: out_word = 8'hFF;
		16'hFBD0: out_word = 8'hFF;
		16'hFBD1: out_word = 8'hFF;
		16'hFBD2: out_word = 8'hFF;
		16'hFBD3: out_word = 8'hFF;
		16'hFBD4: out_word = 8'hFF;
		16'hFBD5: out_word = 8'hFF;
		16'hFBD6: out_word = 8'hFF;
		16'hFBD7: out_word = 8'hFF;
		16'hFBD8: out_word = 8'hFF;
		16'hFBD9: out_word = 8'hFF;
		16'hFBDA: out_word = 8'hFF;
		16'hFBDB: out_word = 8'hFF;
		16'hFBDC: out_word = 8'hFF;
		16'hFBDD: out_word = 8'hFF;
		16'hFBDE: out_word = 8'hFF;
		16'hFBDF: out_word = 8'hFF;
		16'hFBE0: out_word = 8'hFF;
		16'hFBE1: out_word = 8'hFF;
		16'hFBE2: out_word = 8'hFF;
		16'hFBE3: out_word = 8'hFF;
		16'hFBE4: out_word = 8'hFF;
		16'hFBE5: out_word = 8'hFF;
		16'hFBE6: out_word = 8'hFF;
		16'hFBE7: out_word = 8'hFF;
		16'hFBE8: out_word = 8'hFF;
		16'hFBE9: out_word = 8'hFF;
		16'hFBEA: out_word = 8'hFF;
		16'hFBEB: out_word = 8'hFF;
		16'hFBEC: out_word = 8'hFF;
		16'hFBED: out_word = 8'hFF;
		16'hFBEE: out_word = 8'hFF;
		16'hFBEF: out_word = 8'hFF;
		16'hFBF0: out_word = 8'hFF;
		16'hFBF1: out_word = 8'hFF;
		16'hFBF2: out_word = 8'hFF;
		16'hFBF3: out_word = 8'hFF;
		16'hFBF4: out_word = 8'hFF;
		16'hFBF5: out_word = 8'hFF;
		16'hFBF6: out_word = 8'hFF;
		16'hFBF7: out_word = 8'hFF;
		16'hFBF8: out_word = 8'hFF;
		16'hFBF9: out_word = 8'hFF;
		16'hFBFA: out_word = 8'hFF;
		16'hFBFB: out_word = 8'hFF;
		16'hFBFC: out_word = 8'hFF;
		16'hFBFD: out_word = 8'hFF;
		16'hFBFE: out_word = 8'hFF;
		16'hFBFF: out_word = 8'hFF;
		16'hFC00: out_word = 8'hFF;
		16'hFC01: out_word = 8'hFF;
		16'hFC02: out_word = 8'hFF;
		16'hFC03: out_word = 8'hFF;
		16'hFC04: out_word = 8'hFF;
		16'hFC05: out_word = 8'hFF;
		16'hFC06: out_word = 8'hFF;
		16'hFC07: out_word = 8'hFF;
		16'hFC08: out_word = 8'hFF;
		16'hFC09: out_word = 8'hFF;
		16'hFC0A: out_word = 8'hFF;
		16'hFC0B: out_word = 8'hFF;
		16'hFC0C: out_word = 8'hFF;
		16'hFC0D: out_word = 8'hFF;
		16'hFC0E: out_word = 8'hFF;
		16'hFC0F: out_word = 8'hFF;
		16'hFC10: out_word = 8'hFF;
		16'hFC11: out_word = 8'hFF;
		16'hFC12: out_word = 8'hFF;
		16'hFC13: out_word = 8'hFF;
		16'hFC14: out_word = 8'hFF;
		16'hFC15: out_word = 8'hFF;
		16'hFC16: out_word = 8'hFF;
		16'hFC17: out_word = 8'hFF;
		16'hFC18: out_word = 8'hFF;
		16'hFC19: out_word = 8'hFF;
		16'hFC1A: out_word = 8'hFF;
		16'hFC1B: out_word = 8'hFF;
		16'hFC1C: out_word = 8'hFF;
		16'hFC1D: out_word = 8'hFF;
		16'hFC1E: out_word = 8'hFF;
		16'hFC1F: out_word = 8'hFF;
		16'hFC20: out_word = 8'hFF;
		16'hFC21: out_word = 8'hFF;
		16'hFC22: out_word = 8'hFF;
		16'hFC23: out_word = 8'hFF;
		16'hFC24: out_word = 8'hFF;
		16'hFC25: out_word = 8'hFF;
		16'hFC26: out_word = 8'hFF;
		16'hFC27: out_word = 8'hFF;
		16'hFC28: out_word = 8'hFF;
		16'hFC29: out_word = 8'hFF;
		16'hFC2A: out_word = 8'hFF;
		16'hFC2B: out_word = 8'hFF;
		16'hFC2C: out_word = 8'hFF;
		16'hFC2D: out_word = 8'hFF;
		16'hFC2E: out_word = 8'hFF;
		16'hFC2F: out_word = 8'hFF;
		16'hFC30: out_word = 8'hFF;
		16'hFC31: out_word = 8'hFF;
		16'hFC32: out_word = 8'hFF;
		16'hFC33: out_word = 8'hFF;
		16'hFC34: out_word = 8'hFF;
		16'hFC35: out_word = 8'hFF;
		16'hFC36: out_word = 8'hFF;
		16'hFC37: out_word = 8'hFF;
		16'hFC38: out_word = 8'hFF;
		16'hFC39: out_word = 8'hFF;
		16'hFC3A: out_word = 8'hFF;
		16'hFC3B: out_word = 8'hFF;
		16'hFC3C: out_word = 8'hFF;
		16'hFC3D: out_word = 8'hFF;
		16'hFC3E: out_word = 8'hFF;
		16'hFC3F: out_word = 8'hFF;
		16'hFC40: out_word = 8'hFF;
		16'hFC41: out_word = 8'hFF;
		16'hFC42: out_word = 8'hFF;
		16'hFC43: out_word = 8'hFF;
		16'hFC44: out_word = 8'hFF;
		16'hFC45: out_word = 8'hFF;
		16'hFC46: out_word = 8'hFF;
		16'hFC47: out_word = 8'hFF;
		16'hFC48: out_word = 8'hFF;
		16'hFC49: out_word = 8'hFF;
		16'hFC4A: out_word = 8'hFF;
		16'hFC4B: out_word = 8'hFF;
		16'hFC4C: out_word = 8'hFF;
		16'hFC4D: out_word = 8'hFF;
		16'hFC4E: out_word = 8'hFF;
		16'hFC4F: out_word = 8'hFF;
		16'hFC50: out_word = 8'hFF;
		16'hFC51: out_word = 8'hFF;
		16'hFC52: out_word = 8'hFF;
		16'hFC53: out_word = 8'hFF;
		16'hFC54: out_word = 8'hFF;
		16'hFC55: out_word = 8'hFF;
		16'hFC56: out_word = 8'hFF;
		16'hFC57: out_word = 8'hFF;
		16'hFC58: out_word = 8'hFF;
		16'hFC59: out_word = 8'hFF;
		16'hFC5A: out_word = 8'hFF;
		16'hFC5B: out_word = 8'hFF;
		16'hFC5C: out_word = 8'hFF;
		16'hFC5D: out_word = 8'hFF;
		16'hFC5E: out_word = 8'hFF;
		16'hFC5F: out_word = 8'hFF;
		16'hFC60: out_word = 8'hFF;
		16'hFC61: out_word = 8'hFF;
		16'hFC62: out_word = 8'hFF;
		16'hFC63: out_word = 8'hFF;
		16'hFC64: out_word = 8'hFF;
		16'hFC65: out_word = 8'hFF;
		16'hFC66: out_word = 8'hFF;
		16'hFC67: out_word = 8'hFF;
		16'hFC68: out_word = 8'hFF;
		16'hFC69: out_word = 8'hFF;
		16'hFC6A: out_word = 8'hFF;
		16'hFC6B: out_word = 8'hFF;
		16'hFC6C: out_word = 8'hFF;
		16'hFC6D: out_word = 8'hFF;
		16'hFC6E: out_word = 8'hFF;
		16'hFC6F: out_word = 8'hFF;
		16'hFC70: out_word = 8'hFF;
		16'hFC71: out_word = 8'hFF;
		16'hFC72: out_word = 8'hFF;
		16'hFC73: out_word = 8'hFF;
		16'hFC74: out_word = 8'hFF;
		16'hFC75: out_word = 8'hFF;
		16'hFC76: out_word = 8'hFF;
		16'hFC77: out_word = 8'hFF;
		16'hFC78: out_word = 8'hFF;
		16'hFC79: out_word = 8'hFF;
		16'hFC7A: out_word = 8'hFF;
		16'hFC7B: out_word = 8'hFF;
		16'hFC7C: out_word = 8'hFF;
		16'hFC7D: out_word = 8'hFF;
		16'hFC7E: out_word = 8'hFF;
		16'hFC7F: out_word = 8'hFF;
		16'hFC80: out_word = 8'hFF;
		16'hFC81: out_word = 8'hFF;
		16'hFC82: out_word = 8'hFF;
		16'hFC83: out_word = 8'hFF;
		16'hFC84: out_word = 8'hFF;
		16'hFC85: out_word = 8'hFF;
		16'hFC86: out_word = 8'hFF;
		16'hFC87: out_word = 8'hFF;
		16'hFC88: out_word = 8'hFF;
		16'hFC89: out_word = 8'hFF;
		16'hFC8A: out_word = 8'hFF;
		16'hFC8B: out_word = 8'hFF;
		16'hFC8C: out_word = 8'hFF;
		16'hFC8D: out_word = 8'hFF;
		16'hFC8E: out_word = 8'hFF;
		16'hFC8F: out_word = 8'hFF;
		16'hFC90: out_word = 8'hFF;
		16'hFC91: out_word = 8'hFF;
		16'hFC92: out_word = 8'hFF;
		16'hFC93: out_word = 8'hFF;
		16'hFC94: out_word = 8'hFF;
		16'hFC95: out_word = 8'hFF;
		16'hFC96: out_word = 8'hFF;
		16'hFC97: out_word = 8'hFF;
		16'hFC98: out_word = 8'hFF;
		16'hFC99: out_word = 8'hFF;
		16'hFC9A: out_word = 8'hFF;
		16'hFC9B: out_word = 8'hFF;
		16'hFC9C: out_word = 8'hFF;
		16'hFC9D: out_word = 8'hFF;
		16'hFC9E: out_word = 8'hFF;
		16'hFC9F: out_word = 8'hFF;
		16'hFCA0: out_word = 8'hFF;
		16'hFCA1: out_word = 8'hFF;
		16'hFCA2: out_word = 8'hFF;
		16'hFCA3: out_word = 8'hFF;
		16'hFCA4: out_word = 8'hFF;
		16'hFCA5: out_word = 8'hFF;
		16'hFCA6: out_word = 8'hFF;
		16'hFCA7: out_word = 8'hFF;
		16'hFCA8: out_word = 8'hFF;
		16'hFCA9: out_word = 8'hFF;
		16'hFCAA: out_word = 8'hFF;
		16'hFCAB: out_word = 8'hFF;
		16'hFCAC: out_word = 8'hFF;
		16'hFCAD: out_word = 8'hFF;
		16'hFCAE: out_word = 8'hFF;
		16'hFCAF: out_word = 8'hFF;
		16'hFCB0: out_word = 8'hFF;
		16'hFCB1: out_word = 8'hFF;
		16'hFCB2: out_word = 8'hFF;
		16'hFCB3: out_word = 8'hFF;
		16'hFCB4: out_word = 8'hFF;
		16'hFCB5: out_word = 8'hFF;
		16'hFCB6: out_word = 8'hFF;
		16'hFCB7: out_word = 8'hFF;
		16'hFCB8: out_word = 8'hFF;
		16'hFCB9: out_word = 8'hFF;
		16'hFCBA: out_word = 8'hFF;
		16'hFCBB: out_word = 8'hFF;
		16'hFCBC: out_word = 8'hFF;
		16'hFCBD: out_word = 8'hFF;
		16'hFCBE: out_word = 8'hFF;
		16'hFCBF: out_word = 8'hFF;
		16'hFCC0: out_word = 8'hFF;
		16'hFCC1: out_word = 8'hFF;
		16'hFCC2: out_word = 8'hFF;
		16'hFCC3: out_word = 8'hFF;
		16'hFCC4: out_word = 8'hFF;
		16'hFCC5: out_word = 8'hFF;
		16'hFCC6: out_word = 8'hFF;
		16'hFCC7: out_word = 8'hFF;
		16'hFCC8: out_word = 8'hFF;
		16'hFCC9: out_word = 8'hFF;
		16'hFCCA: out_word = 8'hFF;
		16'hFCCB: out_word = 8'hFF;
		16'hFCCC: out_word = 8'hFF;
		16'hFCCD: out_word = 8'hFF;
		16'hFCCE: out_word = 8'hFF;
		16'hFCCF: out_word = 8'hFF;
		16'hFCD0: out_word = 8'hFF;
		16'hFCD1: out_word = 8'hFF;
		16'hFCD2: out_word = 8'hFF;
		16'hFCD3: out_word = 8'hFF;
		16'hFCD4: out_word = 8'hFF;
		16'hFCD5: out_word = 8'hFF;
		16'hFCD6: out_word = 8'hFF;
		16'hFCD7: out_word = 8'hFF;
		16'hFCD8: out_word = 8'hFF;
		16'hFCD9: out_word = 8'hFF;
		16'hFCDA: out_word = 8'hFF;
		16'hFCDB: out_word = 8'hFF;
		16'hFCDC: out_word = 8'hFF;
		16'hFCDD: out_word = 8'hFF;
		16'hFCDE: out_word = 8'hFF;
		16'hFCDF: out_word = 8'hFF;
		16'hFCE0: out_word = 8'hFF;
		16'hFCE1: out_word = 8'hFF;
		16'hFCE2: out_word = 8'hFF;
		16'hFCE3: out_word = 8'hFF;
		16'hFCE4: out_word = 8'hFF;
		16'hFCE5: out_word = 8'hFF;
		16'hFCE6: out_word = 8'hFF;
		16'hFCE7: out_word = 8'hFF;
		16'hFCE8: out_word = 8'hFF;
		16'hFCE9: out_word = 8'hFF;
		16'hFCEA: out_word = 8'hFF;
		16'hFCEB: out_word = 8'hFF;
		16'hFCEC: out_word = 8'hFF;
		16'hFCED: out_word = 8'hFF;
		16'hFCEE: out_word = 8'hFF;
		16'hFCEF: out_word = 8'hFF;
		16'hFCF0: out_word = 8'hFF;
		16'hFCF1: out_word = 8'hFF;
		16'hFCF2: out_word = 8'hFF;
		16'hFCF3: out_word = 8'hFF;
		16'hFCF4: out_word = 8'hFF;
		16'hFCF5: out_word = 8'hFF;
		16'hFCF6: out_word = 8'hFF;
		16'hFCF7: out_word = 8'hFF;
		16'hFCF8: out_word = 8'hFF;
		16'hFCF9: out_word = 8'hFF;
		16'hFCFA: out_word = 8'hFF;
		16'hFCFB: out_word = 8'hFF;
		16'hFCFC: out_word = 8'hFF;
		16'hFCFD: out_word = 8'hFF;
		16'hFCFE: out_word = 8'hFF;
		16'hFCFF: out_word = 8'hFF;
		16'hFD00: out_word = 8'hFF;
		16'hFD01: out_word = 8'hFF;
		16'hFD02: out_word = 8'hFF;
		16'hFD03: out_word = 8'hFF;
		16'hFD04: out_word = 8'hFF;
		16'hFD05: out_word = 8'hFF;
		16'hFD06: out_word = 8'hFF;
		16'hFD07: out_word = 8'hFF;
		16'hFD08: out_word = 8'hFF;
		16'hFD09: out_word = 8'hFF;
		16'hFD0A: out_word = 8'hFF;
		16'hFD0B: out_word = 8'hFF;
		16'hFD0C: out_word = 8'hFF;
		16'hFD0D: out_word = 8'hFF;
		16'hFD0E: out_word = 8'hFF;
		16'hFD0F: out_word = 8'hFF;
		16'hFD10: out_word = 8'hFF;
		16'hFD11: out_word = 8'hFF;
		16'hFD12: out_word = 8'hFF;
		16'hFD13: out_word = 8'hFF;
		16'hFD14: out_word = 8'hFF;
		16'hFD15: out_word = 8'hFF;
		16'hFD16: out_word = 8'hFF;
		16'hFD17: out_word = 8'hFF;
		16'hFD18: out_word = 8'hFF;
		16'hFD19: out_word = 8'hFF;
		16'hFD1A: out_word = 8'hFF;
		16'hFD1B: out_word = 8'hFF;
		16'hFD1C: out_word = 8'hFF;
		16'hFD1D: out_word = 8'hFF;
		16'hFD1E: out_word = 8'hFF;
		16'hFD1F: out_word = 8'hFF;
		16'hFD20: out_word = 8'hFF;
		16'hFD21: out_word = 8'hFF;
		16'hFD22: out_word = 8'hFF;
		16'hFD23: out_word = 8'hFF;
		16'hFD24: out_word = 8'hFF;
		16'hFD25: out_word = 8'hFF;
		16'hFD26: out_word = 8'hFF;
		16'hFD27: out_word = 8'hFF;
		16'hFD28: out_word = 8'hFF;
		16'hFD29: out_word = 8'hFF;
		16'hFD2A: out_word = 8'hFF;
		16'hFD2B: out_word = 8'hFF;
		16'hFD2C: out_word = 8'hFF;
		16'hFD2D: out_word = 8'hFF;
		16'hFD2E: out_word = 8'hFF;
		16'hFD2F: out_word = 8'h00;
		16'hFD30: out_word = 8'hC9;
		16'hFD31: out_word = 8'h01;
		16'hFD32: out_word = 8'hFD;
		16'hFD33: out_word = 8'h7F;
		16'hFD34: out_word = 8'h3E;
		16'hFD35: out_word = 8'h10;
		16'hFD36: out_word = 8'hED;
		16'hFD37: out_word = 8'h79;
		16'hFD38: out_word = 8'hFB;
		16'hFD39: out_word = 8'h21;
		16'hFD3A: out_word = 8'hBF;
		16'hFD3B: out_word = 8'h80;
		16'hFD3C: out_word = 8'h11;
		16'hFD3D: out_word = 8'hC0;
		16'hFD3E: out_word = 8'h80;
		16'hFD3F: out_word = 8'h7B;
		16'hFD40: out_word = 8'h87;
		16'hFD41: out_word = 8'h87;
		16'hFD42: out_word = 8'hD9;
		16'hFD43: out_word = 8'h16;
		16'hFD44: out_word = 8'h00;
		16'hFD45: out_word = 8'h5F;
		16'hFD46: out_word = 8'h62;
		16'hFD47: out_word = 8'h6A;
		16'hFD48: out_word = 8'h19;
		16'hFD49: out_word = 8'h3D;
		16'hFD4A: out_word = 8'h20;
		16'hFD4B: out_word = 8'hFC;
		16'hFD4C: out_word = 8'h7C;
		16'hFD4D: out_word = 8'h37;
		16'hFD4E: out_word = 8'h1F;
		16'hFD4F: out_word = 8'hD9;
		16'hFD50: out_word = 8'h12;
		16'hFD51: out_word = 8'h77;
		16'hFD52: out_word = 8'hCB;
		16'hFD53: out_word = 8'hBD;
		16'hFD54: out_word = 8'hCB;
		16'hFD55: out_word = 8'hBB;
		16'hFD56: out_word = 8'h2F;
		16'hFD57: out_word = 8'h12;
		16'hFD58: out_word = 8'h77;
		16'hFD59: out_word = 8'hCB;
		16'hFD5A: out_word = 8'hFD;
		16'hFD5B: out_word = 8'hCB;
		16'hFD5C: out_word = 8'hFB;
		16'hFD5D: out_word = 8'h2D;
		16'hFD5E: out_word = 8'h1C;
		16'hFD5F: out_word = 8'h20;
		16'hFD60: out_word = 8'hDE;
		16'hFD61: out_word = 8'h24;
		16'hFD62: out_word = 8'h36;
		16'hFD63: out_word = 8'hB0;
		16'hFD64: out_word = 8'h2C;
		16'hFD65: out_word = 8'h73;
		16'hFD66: out_word = 8'h23;
		16'hFD67: out_word = 8'h7C;
		16'hFD68: out_word = 8'hFE;
		16'hFD69: out_word = 8'h58;
		16'hFD6A: out_word = 8'h20;
		16'hFD6B: out_word = 8'hF9;
		16'hFD6C: out_word = 8'h76;
		16'hFD6D: out_word = 8'h11;
		16'hFD6E: out_word = 8'h04;
		16'hFD6F: out_word = 8'h0D;
		16'hFD70: out_word = 8'h3E;
		16'hFD71: out_word = 8'h01;
		16'hFD72: out_word = 8'h3D;
		16'hFD73: out_word = 8'h20;
		16'hFD74: out_word = 8'h69;
		16'hFD75: out_word = 8'hD3;
		16'hFD76: out_word = 8'hFE;
		16'hFD77: out_word = 8'h21;
		16'hFD78: out_word = 8'hD8;
		16'hFD79: out_word = 8'h61;
		16'hFD7A: out_word = 8'h06;
		16'hFD7B: out_word = 8'h08;
		16'hFD7C: out_word = 8'h3E;
		16'hFD7D: out_word = 8'h41;
		16'hFD7E: out_word = 8'hCD;
		16'hFD7F: out_word = 8'hEE;
		16'hFD80: out_word = 8'h61;
		16'hFD81: out_word = 8'h07;
		16'hFD82: out_word = 8'hCD;
		16'hFD83: out_word = 8'hEE;
		16'hFD84: out_word = 8'h61;
		16'hFD85: out_word = 8'h07;
		16'hFD86: out_word = 8'h07;
		16'hFD87: out_word = 8'h32;
		16'hFD88: out_word = 8'hEB;
		16'hFD89: out_word = 8'h61;
		16'hFD8A: out_word = 8'hD6;
		16'hFD8B: out_word = 8'h38;
		16'hFD8C: out_word = 8'h28;
		16'hFD8D: out_word = 8'h02;
		16'hFD8E: out_word = 8'h3E;
		16'hFD8F: out_word = 8'h10;
		16'hFD90: out_word = 8'h32;
		16'hFD91: out_word = 8'hE8;
		16'hFD92: out_word = 8'h61;
		16'hFD93: out_word = 8'h2B;
		16'hFD94: out_word = 8'hCB;
		16'hFD95: out_word = 8'h0E;
		16'hFD96: out_word = 8'h30;
		16'hFD97: out_word = 8'h0D;
		16'hFD98: out_word = 8'hD9;
		16'hFD99: out_word = 8'h3E;
		16'hFD9A: out_word = 8'h10;
		16'hFD9B: out_word = 8'h32;
		16'hFD9C: out_word = 8'hE9;
		16'hFD9D: out_word = 8'h61;
		16'hFD9E: out_word = 8'h21;
		16'hFD9F: out_word = 8'hBB;
		16'hFDA0: out_word = 8'h81;
		16'hFDA1: out_word = 8'hCD;
		16'hFDA2: out_word = 8'hBD;
		16'hFDA3: out_word = 8'h61;
		16'hFDA4: out_word = 8'hD9;
		16'hFDA5: out_word = 8'h21;
		16'hFDA6: out_word = 8'hFF;
		16'hFDA7: out_word = 8'hFF;
		16'hFDA8: out_word = 8'h23;
		16'hFDA9: out_word = 8'h22;
		16'hFDAA: out_word = 8'h6D;
		16'hFDAB: out_word = 8'h60;
		16'hFDAC: out_word = 8'h29;
		16'hFDAD: out_word = 8'h7D;
		16'hFDAE: out_word = 8'hB7;
		16'hFDAF: out_word = 8'h20;
		16'hFDB0: out_word = 8'h01;
		16'hFDB1: out_word = 8'h14;
		16'hFDB2: out_word = 8'h7C;
		16'hFDB3: out_word = 8'hE6;
		16'hFDB4: out_word = 8'h03;
		16'hFDB5: out_word = 8'h28;
		16'hFDB6: out_word = 8'h25;
		16'hFDB7: out_word = 8'h06;
		16'hFDB8: out_word = 8'h01;
		16'hFDB9: out_word = 8'h3D;
		16'hFDBA: out_word = 8'h20;
		16'hFDBB: out_word = 8'h02;
		16'hFDBC: out_word = 8'h06;
		16'hFDBD: out_word = 8'h04;
		16'hFDBE: out_word = 8'hAF;
		16'hFDBF: out_word = 8'h21;
		16'hFDC0: out_word = 8'hE0;
		16'hFDC1: out_word = 8'h61;
		16'hFDC2: out_word = 8'hCD;
		16'hFDC3: out_word = 8'hEE;
		16'hFDC4: out_word = 8'h61;
		16'hFDC5: out_word = 8'h87;
		16'hFDC6: out_word = 8'h28;
		16'hFDC7: out_word = 8'h14;
		16'hFDC8: out_word = 8'h32;
		16'hFDC9: out_word = 8'hE5;
		16'hFDCA: out_word = 8'h61;
		16'hFDCB: out_word = 8'h3E;
		16'hFDCC: out_word = 8'h10;
		16'hFDCD: out_word = 8'h32;
		16'hFDCE: out_word = 8'hEA;
		16'hFDCF: out_word = 8'h61;
		16'hFDD0: out_word = 8'h1E;
		16'hFDD1: out_word = 8'h47;
		16'hFDD2: out_word = 8'hD9;
		16'hFDD3: out_word = 8'h3E;
		16'hFDD4: out_word = 8'h30;
		16'hFDD5: out_word = 8'h21;
		16'hFDD6: out_word = 8'h8B;
		16'hFDD7: out_word = 8'h81;
		16'hFDD8: out_word = 8'hCD;
		16'hFDD9: out_word = 8'hBD;
		16'hFDDA: out_word = 8'h61;
		16'hFDDB: out_word = 8'hD9;
		16'hFDDC: out_word = 8'h3E;
		16'hFDDD: out_word = 8'h05;
		16'hFDDE: out_word = 8'h32;
		16'hFDDF: out_word = 8'h38;
		16'hFDE0: out_word = 8'h60;
		16'hFDE1: out_word = 8'h21;
		16'hFDE2: out_word = 8'hE9;
		16'hFDE3: out_word = 8'h61;
		16'hFDE4: out_word = 8'h0F;
		16'hFDE5: out_word = 8'hD4;
		16'hFDE6: out_word = 8'hD2;
		16'hFDE7: out_word = 8'h61;
		16'hFDE8: out_word = 8'h23;
		16'hFDE9: out_word = 8'hCD;
		16'hFDEA: out_word = 8'hD2;
		16'hFDEB: out_word = 8'h61;
		16'hFDEC: out_word = 8'h7E;
		16'hFDED: out_word = 8'h0F;
		16'hFDEE: out_word = 8'h0F;
		16'hFDEF: out_word = 8'hE6;
		16'hFDF0: out_word = 8'h03;
		16'hFDF1: out_word = 8'h3C;
		16'hFDF2: out_word = 8'h08;
		16'hFDF3: out_word = 8'h21;
		16'hFDF4: out_word = 8'hE5;
		16'hFDF5: out_word = 8'h61;
		16'hFDF6: out_word = 8'h34;
		16'hFDF7: out_word = 8'h2B;
		16'hFDF8: out_word = 8'h3E;
		16'hFDF9: out_word = 8'h04;
		16'hFDFA: out_word = 8'h01;
		16'hFDFB: out_word = 8'hFD;
		16'hFDFC: out_word = 8'hFF;
		16'hFDFD: out_word = 8'hED;
		16'hFDFE: out_word = 8'h79;
		16'hFDFF: out_word = 8'h06;
		16'hFE00: out_word = 8'hBF;
		16'hFE01: out_word = 8'hED;
		16'hFE02: out_word = 8'hA3;
		16'hFE03: out_word = 8'h3C;
		16'hFE04: out_word = 8'hBA;
		16'hFE05: out_word = 8'h20;
		16'hFE06: out_word = 8'hF3;
		16'hFE07: out_word = 8'h21;
		16'hFE08: out_word = 8'h00;
		16'hFE09: out_word = 8'h58;
		16'hFE0A: out_word = 8'h73;
		16'hFE0B: out_word = 8'h11;
		16'hFE0C: out_word = 8'h01;
		16'hFE0D: out_word = 8'h58;
		16'hFE0E: out_word = 8'h01;
		16'hFE0F: out_word = 8'hFF;
		16'hFE10: out_word = 8'h02;
		16'hFE11: out_word = 8'hED;
		16'hFE12: out_word = 8'hB0;
		16'hFE13: out_word = 8'h08;
		16'hFE14: out_word = 8'h4F;
		16'hFE15: out_word = 8'h06;
		16'hFE16: out_word = 8'h06;
		16'hFE17: out_word = 8'h21;
		16'hFE18: out_word = 8'h7F;
		16'hFE19: out_word = 8'h81;
		16'hFE1A: out_word = 8'hC5;
		16'hFE1B: out_word = 8'h7E;
		16'hFE1C: out_word = 8'h2C;
		16'hFE1D: out_word = 8'hE5;
		16'hFE1E: out_word = 8'h07;
		16'hFE1F: out_word = 8'h30;
		16'hFE20: out_word = 8'h59;
		16'hFE21: out_word = 8'h07;
		16'hFE22: out_word = 8'h35;
		16'hFE23: out_word = 8'h20;
		16'hFE24: out_word = 8'h06;
		16'hFE25: out_word = 8'h30;
		16'hFE26: out_word = 8'h04;
		16'hFE27: out_word = 8'hAF;
		16'hFE28: out_word = 8'h2D;
		16'hFE29: out_word = 8'h77;
		16'hFE2A: out_word = 8'h2C;
		16'hFE2B: out_word = 8'h2C;
		16'hFE2C: out_word = 8'h11;
		16'hFE2D: out_word = 8'h00;
		16'hFE2E: out_word = 8'h00;
		16'hFE2F: out_word = 8'h01;
		16'hFE30: out_word = 8'hA6;
		16'hFE31: out_word = 8'h61;
		16'hFE32: out_word = 8'hCD;
		16'hFE33: out_word = 8'h90;
		16'hFE34: out_word = 8'h61;
		16'hFE35: out_word = 8'h01;
		16'hFE36: out_word = 8'h79;
		16'hFE37: out_word = 8'h61;
		16'hFE38: out_word = 8'hCD;
		16'hFE39: out_word = 8'h90;
		16'hFE3A: out_word = 8'h61;
		16'hFE3B: out_word = 8'h08;
		16'hFE3C: out_word = 8'hCD;
		16'hFE3D: out_word = 8'h8D;
		16'hFE3E: out_word = 8'h61;
		16'hFE3F: out_word = 8'hD5;
		16'hFE40: out_word = 8'h7A;
		16'hFE41: out_word = 8'hCD;
		16'hFE42: out_word = 8'hB3;
		16'hFE43: out_word = 8'h61;
		16'hFE44: out_word = 8'hCD;
		16'hFE45: out_word = 8'h8D;
		16'hFE46: out_word = 8'h61;
		16'hFE47: out_word = 8'hF1;
		16'hFE48: out_word = 8'hD5;
		16'hFE49: out_word = 8'hC6;
		16'hFE4A: out_word = 8'h40;
		16'hFE4B: out_word = 8'hCD;
		16'hFE4C: out_word = 8'hB3;
		16'hFE4D: out_word = 8'h61;
		16'hFE4E: out_word = 8'h01;
		16'hFE4F: out_word = 8'h83;
		16'hFE50: out_word = 8'h61;
		16'hFE51: out_word = 8'hCD;
		16'hFE52: out_word = 8'h90;
		16'hFE53: out_word = 8'h61;
		16'hFE54: out_word = 8'hC1;
		16'hFE55: out_word = 8'hCD;
		16'hFE56: out_word = 8'h4F;
		16'hFE57: out_word = 8'h61;
		16'hFE58: out_word = 8'h08;
		16'hFE59: out_word = 8'h07;
		16'hFE5A: out_word = 8'h30;
		16'hFE5B: out_word = 8'h1E;
		16'hFE5C: out_word = 8'hCD;
		16'hFE5D: out_word = 8'hA7;
		16'hFE5E: out_word = 8'h61;
		16'hFE5F: out_word = 8'hFE;
		16'hFE60: out_word = 8'hF0;
		16'hFE61: out_word = 8'h38;
		16'hFE62: out_word = 8'h17;
		16'hFE63: out_word = 8'h06;
		16'hFE64: out_word = 8'h04;
		16'hFE65: out_word = 8'h21;
		16'hFE66: out_word = 8'h8B;
		16'hFE67: out_word = 8'h81;
		16'hFE68: out_word = 8'h11;
		16'hFE69: out_word = 8'h0C;
		16'hFE6A: out_word = 8'h00;
		16'hFE6B: out_word = 8'hCB;
		16'hFE6C: out_word = 8'h7E;
		16'hFE6D: out_word = 8'h20;
		16'hFE6E: out_word = 8'h08;
		16'hFE6F: out_word = 8'hD1;
		16'hFE70: out_word = 8'hD5;
		16'hFE71: out_word = 8'h1A;
		16'hFE72: out_word = 8'h1D;
		16'hFE73: out_word = 8'hCD;
		16'hFE74: out_word = 8'hC0;
		16'hFE75: out_word = 8'h61;
		16'hFE76: out_word = 8'h04;
		16'hFE77: out_word = 8'h19;
		16'hFE78: out_word = 8'h10;
		16'hFE79: out_word = 8'hF1;
		16'hFE7A: out_word = 8'hE1;
		16'hFE7B: out_word = 8'h01;
		16'hFE7C: out_word = 8'h0B;
		16'hFE7D: out_word = 8'h00;
		16'hFE7E: out_word = 8'h09;
		16'hFE7F: out_word = 8'hC1;
		16'hFE80: out_word = 8'h10;
		16'hFE81: out_word = 8'h98;
		16'hFE82: out_word = 8'h0D;
		16'hFE83: out_word = 8'h20;
		16'hFE84: out_word = 8'h90;
		16'hFE85: out_word = 8'hC3;
		16'hFE86: out_word = 8'h33;
		16'hFE87: out_word = 8'h60;
		16'hFE88: out_word = 8'h21;
		16'hFE89: out_word = 8'h00;
		16'hFE8A: out_word = 8'hC0;
		16'hFE8B: out_word = 8'h58;
		16'hFE8C: out_word = 8'h4E;
		16'hFE8D: out_word = 8'h73;
		16'hFE8E: out_word = 8'h2C;
		16'hFE8F: out_word = 8'h7E;
		16'hFE90: out_word = 8'h72;
		16'hFE91: out_word = 8'h23;
		16'hFE92: out_word = 8'hCB;
		16'hFE93: out_word = 8'h9C;
		16'hFE94: out_word = 8'h22;
		16'hFE95: out_word = 8'h50;
		16'hFE96: out_word = 8'h61;
		16'hFE97: out_word = 8'h21;
		16'hFE98: out_word = 8'h2F;
		16'hFE99: out_word = 8'hA6;
		16'hFE9A: out_word = 8'hCD;
		16'hFE9B: out_word = 8'h69;
		16'hFE9C: out_word = 8'h61;
		16'hFE9D: out_word = 8'h7A;
		16'hFE9E: out_word = 8'h4B;
		16'hFE9F: out_word = 8'h21;
		16'hFEA0: out_word = 8'h00;
		16'hFEA1: out_word = 8'hB6;
		16'hFEA2: out_word = 8'h22;
		16'hFEA3: out_word = 8'h76;
		16'hFEA4: out_word = 8'h61;
		16'hFEA5: out_word = 8'hCD;
		16'hFEA6: out_word = 8'hB0;
		16'hFEA7: out_word = 8'h22;
		16'hFEA8: out_word = 8'h3C;
		16'hFEA9: out_word = 8'h47;
		16'hFEAA: out_word = 8'h3E;
		16'hFEAB: out_word = 8'h01;
		16'hFEAC: out_word = 8'h0F;
		16'hFEAD: out_word = 8'h10;
		16'hFEAE: out_word = 8'hFD;
		16'hFEAF: out_word = 8'h2F;
		16'hFEB0: out_word = 8'hA6;
		16'hFEB1: out_word = 8'h77;
		16'hFEB2: out_word = 8'hD0;
		16'hFEB3: out_word = 8'h7A;
		16'hFEB4: out_word = 8'h07;
		16'hFEB5: out_word = 8'h9F;
		16'hFEB6: out_word = 8'hAA;
		16'hFEB7: out_word = 8'hE6;
		16'hFEB8: out_word = 8'hFE;
		16'hFEB9: out_word = 8'hAA;
		16'hFEBA: out_word = 8'h57;
		16'hFEBB: out_word = 8'hC9;
		16'hFEBC: out_word = 8'h7A;
		16'hFEBD: out_word = 8'hFE;
		16'hFEBE: out_word = 8'hC0;
		16'hFEBF: out_word = 8'hD8;
		16'hFEC0: out_word = 8'h0F;
		16'hFEC1: out_word = 8'h9F;
		16'hFEC2: out_word = 8'hE6;
		16'hFEC3: out_word = 8'hBF;
		16'hFEC4: out_word = 8'h57;
		16'hFEC5: out_word = 8'hC9;
		16'hFEC6: out_word = 8'h01;
		16'hFEC7: out_word = 8'hA5;
		16'hFEC8: out_word = 8'h61;
		16'hFEC9: out_word = 8'hED;
		16'hFECA: out_word = 8'h43;
		16'hFECB: out_word = 8'h9E;
		16'hFECC: out_word = 8'h61;
		16'hFECD: out_word = 8'h4E;
		16'hFECE: out_word = 8'h2C;
		16'hFECF: out_word = 8'h46;
		16'hFED0: out_word = 8'h2D;
		16'hFED1: out_word = 8'hEB;
		16'hFED2: out_word = 8'h09;
		16'hFED3: out_word = 8'hEB;
		16'hFED4: out_word = 8'h07;
		16'hFED5: out_word = 8'hF5;
		16'hFED6: out_word = 8'hCD;
		16'hFED7: out_word = 8'hA5;
		16'hFED8: out_word = 8'h61;
		16'hFED9: out_word = 8'hF1;
		16'hFEDA: out_word = 8'h73;
		16'hFEDB: out_word = 8'h2C;
		16'hFEDC: out_word = 8'h72;
		16'hFEDD: out_word = 8'h2C;
		16'hFEDE: out_word = 8'hC9;
		16'hFEDF: out_word = 8'hD0;
		16'hFEE0: out_word = 8'h11;
		16'hFEE1: out_word = 8'hE0;
		16'hFEE2: out_word = 8'h17;
		16'hFEE3: out_word = 8'h13;
		16'hFEE4: out_word = 8'hCB;
		16'hFEE5: out_word = 8'hAA;
		16'hFEE6: out_word = 8'hED;
		16'hFEE7: out_word = 8'h53;
		16'hFEE8: out_word = 8'hA8;
		16'hFEE9: out_word = 8'h61;
		16'hFEEA: out_word = 8'h18;
		16'hFEEB: out_word = 8'h03;
		16'hFEEC: out_word = 8'h16;
		16'hFEED: out_word = 8'h80;
		16'hFEEE: out_word = 8'h5F;
		16'hFEEF: out_word = 8'h1A;
		16'hFEF0: out_word = 8'h07;
		16'hFEF1: out_word = 8'h5F;
		16'hFEF2: out_word = 8'h9F;
		16'hFEF3: out_word = 8'h57;
		16'hFEF4: out_word = 8'h7B;
		16'hFEF5: out_word = 8'hC9;
		16'hFEF6: out_word = 8'h11;
		16'hFEF7: out_word = 8'h7F;
		16'hFEF8: out_word = 8'h81;
		16'hFEF9: out_word = 8'hE5;
		16'hFEFA: out_word = 8'hEB;
		16'hFEFB: out_word = 8'h01;
		16'hFEFC: out_word = 8'h0C;
		16'hFEFD: out_word = 8'h00;
		16'hFEFE: out_word = 8'hED;
		16'hFEFF: out_word = 8'hB0;
		16'hFF00: out_word = 8'hE1;
		16'hFF01: out_word = 8'h36;
		16'hFF02: out_word = 8'hC8;
		16'hFF03: out_word = 8'h2C;
		16'hFF04: out_word = 8'h77;
		16'hFF05: out_word = 8'h2C;
		16'hFF06: out_word = 8'hCD;
		16'hFF07: out_word = 8'hA7;
		16'hFF08: out_word = 8'h61;
		16'hFF09: out_word = 8'h18;
		16'hFF0A: out_word = 8'hCF;
		16'hFF0B: out_word = 8'h7E;
		16'hFF0C: out_word = 8'h3D;
		16'hFF0D: out_word = 8'hF8;
		16'hFF0E: out_word = 8'h35;
		16'hFF0F: out_word = 8'hC9;
		16'hFF10: out_word = 8'h44;
		16'hFF11: out_word = 8'h0A;
		16'hFF12: out_word = 8'h66;
		16'hFF13: out_word = 8'hA0;
		16'hFF14: out_word = 8'h00;
		16'hFF15: out_word = 8'hF7;
		16'hFF16: out_word = 8'h77;
		16'hFF17: out_word = 8'hF7;
		16'hFF18: out_word = 8'hFF;
		16'hFF19: out_word = 8'h11;
		16'hFF1A: out_word = 8'h11;
		16'hFF1B: out_word = 8'h14;
		16'hFF1C: out_word = 8'h41;
		16'hFF1D: out_word = 8'hDF;
		16'hFF1E: out_word = 8'h01;
		16'hFF1F: out_word = 8'h00;
		16'hFF20: out_word = 8'h2B;
		16'hFF21: out_word = 8'h00;
		16'hFF22: out_word = 8'h00;
		16'hFF23: out_word = 8'h00;
		16'hFF24: out_word = 8'h00;
		16'hFF25: out_word = 8'h00;
		16'hFF26: out_word = 8'h0E;
		16'hFF27: out_word = 8'hC5;
		16'hFF28: out_word = 8'hE5;
		16'hFF29: out_word = 8'h4E;
		16'hFF2A: out_word = 8'hCB;
		16'hFF2B: out_word = 8'h1E;
		16'hFF2C: out_word = 8'h2C;
		16'hFF2D: out_word = 8'h10;
		16'hFF2E: out_word = 8'hFB;
		16'hFF2F: out_word = 8'hE1;
		16'hFF30: out_word = 8'hF5;
		16'hFF31: out_word = 8'hCB;
		16'hFF32: out_word = 8'h19;
		16'hFF33: out_word = 8'h71;
		16'hFF34: out_word = 8'hF1;
		16'hFF35: out_word = 8'hC1;
		16'hFF36: out_word = 8'h17;
		16'hFF37: out_word = 8'hC9;
		16'hFF38: out_word = 8'h3E;
		16'hFF39: out_word = 8'h80;
		16'hFF3A: out_word = 8'h08;
		16'hFF3B: out_word = 8'hED;
		16'hFF3C: out_word = 8'hA0;
		16'hFF3D: out_word = 8'h01;
		16'hFF3E: out_word = 8'hFF;
		16'hFF3F: out_word = 8'h02;
		16'hFF40: out_word = 8'h08;
		16'hFF41: out_word = 8'h87;
		16'hFF42: out_word = 8'h20;
		16'hFF43: out_word = 8'h03;
		16'hFF44: out_word = 8'h7E;
		16'hFF45: out_word = 8'h23;
		16'hFF46: out_word = 8'h17;
		16'hFF47: out_word = 8'hCB;
		16'hFF48: out_word = 8'h11;
		16'hFF49: out_word = 8'h30;
		16'hFF4A: out_word = 8'hF6;
		16'hFF4B: out_word = 8'h08;
		16'hFF4C: out_word = 8'h10;
		16'hFF4D: out_word = 8'h0F;
		16'hFF4E: out_word = 8'h3E;
		16'hFF4F: out_word = 8'h02;
		16'hFF50: out_word = 8'hCB;
		16'hFF51: out_word = 8'h29;
		16'hFF52: out_word = 8'h38;
		16'hFF53: out_word = 8'h18;
		16'hFF54: out_word = 8'h3C;
		16'hFF55: out_word = 8'h0C;
		16'hFF56: out_word = 8'h28;
		16'hFF57: out_word = 8'h0F;
		16'hFF58: out_word = 8'h01;
		16'hFF59: out_word = 8'h3F;
		16'hFF5A: out_word = 8'h03;
		16'hFF5B: out_word = 8'h18;
		16'hFF5C: out_word = 8'hE3;
		16'hFF5D: out_word = 8'h10;
		16'hFF5E: out_word = 8'h25;
		16'hFF5F: out_word = 8'hCB;
		16'hFF60: out_word = 8'h39;
		16'hFF61: out_word = 8'h38;
		16'hFF62: out_word = 8'hD8;
		16'hFF63: out_word = 8'h04;
		16'hFF64: out_word = 8'h18;
		16'hFF65: out_word = 8'hDA;
		16'hFF66: out_word = 8'h81;
		16'hFF67: out_word = 8'h01;
		16'hFF68: out_word = 8'hFF;
		16'hFF69: out_word = 8'h04;
		16'hFF6A: out_word = 8'h18;
		16'hFF6B: out_word = 8'hD4;
		16'hFF6C: out_word = 8'h0C;
		16'hFF6D: out_word = 8'h20;
		16'hFF6E: out_word = 8'h28;
		16'hFF6F: out_word = 8'h08;
		16'hFF70: out_word = 8'h04;
		16'hFF71: out_word = 8'hCB;
		16'hFF72: out_word = 8'h19;
		16'hFF73: out_word = 8'hD8;
		16'hFF74: out_word = 8'hCB;
		16'hFF75: out_word = 8'h10;
		16'hFF76: out_word = 8'h87;
		16'hFF77: out_word = 8'h20;
		16'hFF78: out_word = 8'h03;
		16'hFF79: out_word = 8'h7E;
		16'hFF7A: out_word = 8'h23;
		16'hFF7B: out_word = 8'h17;
		16'hFF7C: out_word = 8'h30;
		16'hFF7D: out_word = 8'hF3;
		16'hFF7E: out_word = 8'h08;
		16'hFF7F: out_word = 8'h80;
		16'hFF80: out_word = 8'h06;
		16'hFF81: out_word = 8'h06;
		16'hFF82: out_word = 8'h18;
		16'hFF83: out_word = 8'hBC;
		16'hFF84: out_word = 8'h10;
		16'hFF85: out_word = 8'h04;
		16'hFF86: out_word = 8'h3E;
		16'hFF87: out_word = 8'h01;
		16'hFF88: out_word = 8'h18;
		16'hFF89: out_word = 8'h0F;
		16'hFF8A: out_word = 8'h10;
		16'hFF8B: out_word = 8'h08;
		16'hFF8C: out_word = 8'h0C;
		16'hFF8D: out_word = 8'h20;
		16'hFF8E: out_word = 8'h08;
		16'hFF8F: out_word = 8'h01;
		16'hFF90: out_word = 8'h1F;
		16'hFF91: out_word = 8'h05;
		16'hFF92: out_word = 8'h18;
		16'hFF93: out_word = 8'hAC;
		16'hFF94: out_word = 8'h10;
		16'hFF95: out_word = 8'hD0;
		16'hFF96: out_word = 8'h41;
		16'hFF97: out_word = 8'h4E;
		16'hFF98: out_word = 8'h23;
		16'hFF99: out_word = 8'h05;
		16'hFF9A: out_word = 8'hE5;
		16'hFF9B: out_word = 8'h69;
		16'hFF9C: out_word = 8'h60;
		16'hFF9D: out_word = 8'h19;
		16'hFF9E: out_word = 8'h4F;
		16'hFF9F: out_word = 8'h06;
		16'hFFA0: out_word = 8'h00;
		16'hFFA1: out_word = 8'hED;
		16'hFFA2: out_word = 8'hB0;
		16'hFFA3: out_word = 8'hE1;
		16'hFFA4: out_word = 8'h18;
		16'hFFA5: out_word = 8'h97;
		16'hFFA6: out_word = 8'h83;
		16'hFFA7: out_word = 8'h7A;
		16'hFFA8: out_word = 8'h7D;
		16'hFFA9: out_word = 8'hFF;
		16'hFFAA: out_word = 8'h00;
		16'hFFAB: out_word = 8'h7A;
		16'hFFAC: out_word = 8'h7D;
		16'hFFAD: out_word = 8'hFF;
		16'hFFAE: out_word = 8'hF1;
		16'hFFAF: out_word = 8'hE1;
		16'hFFB0: out_word = 8'hD1;
		16'hFFB1: out_word = 8'hC1;
		16'hFFB2: out_word = 8'hC1;
		16'hFFB3: out_word = 8'hB1;
		16'hFFB4: out_word = 8'hA1;
		16'hFFB5: out_word = 8'h91;
		16'hFFB6: out_word = 8'h41;
		16'hFFB7: out_word = 8'h21;
		16'hFFB8: out_word = 8'h31;
		16'hFFB9: out_word = 8'h11;
		16'hFFBA: out_word = 8'h01;
		16'hFFBB: out_word = 8'h01;
		16'hFFBC: out_word = 8'hF1;
		16'hFFBD: out_word = 8'hE1;
		16'hFFBE: out_word = 8'h00;
		16'hFFBF: out_word = 8'h21;
		16'hFFC0: out_word = 8'h42;
		16'hFFC1: out_word = 8'h63;
		16'hFFC2: out_word = 8'h90;
		16'hFFC3: out_word = 8'hB1;
		16'hFFC4: out_word = 8'hD2;
		16'hFFC5: out_word = 8'hF3;
		16'hFFC6: out_word = 8'hE0;
		16'hFFC7: out_word = 8'hE1;
		16'hFFC8: out_word = 8'hE2;
		16'hFFC9: out_word = 8'hE3;
		16'hFFCA: out_word = 8'hF0;
		16'hFFCB: out_word = 8'hF1;
		16'hFFCC: out_word = 8'hF2;
		16'hFFCD: out_word = 8'hF3;
		16'hFFCE: out_word = 8'hFF;
		16'hFFCF: out_word = 8'hFF;
		16'hFFD0: out_word = 8'hFF;
		16'hFFD1: out_word = 8'hFF;
		16'hFFD2: out_word = 8'hFF;
		16'hFFD3: out_word = 8'hFF;
		16'hFFD4: out_word = 8'hFF;
		16'hFFD5: out_word = 8'hFF;
		16'hFFD6: out_word = 8'hFF;
		16'hFFD7: out_word = 8'hFF;
		16'hFFD8: out_word = 8'hFF;
		16'hFFD9: out_word = 8'hFF;
		16'hFFDA: out_word = 8'hFF;
		16'hFFDB: out_word = 8'hFF;
		16'hFFDC: out_word = 8'hFF;
		16'hFFDD: out_word = 8'hFF;
		16'hFFDE: out_word = 8'hFF;
		16'hFFDF: out_word = 8'hFF;
		16'hFFE0: out_word = 8'hFF;
		16'hFFE1: out_word = 8'hFF;
		16'hFFE2: out_word = 8'hFF;
		16'hFFE3: out_word = 8'hFF;
		16'hFFE4: out_word = 8'hFF;
		16'hFFE5: out_word = 8'hFF;
		16'hFFE6: out_word = 8'hFF;
		16'hFFE7: out_word = 8'hFF;
		16'hFFE8: out_word = 8'hFF;
		16'hFFE9: out_word = 8'hFF;
		16'hFFEA: out_word = 8'hFF;
		16'hFFEB: out_word = 8'hFF;
		16'hFFEC: out_word = 8'hFF;
		16'hFFED: out_word = 8'hFF;
		16'hFFEE: out_word = 8'hFF;
		16'hFFEF: out_word = 8'hFF;
		16'hFFF0: out_word = 8'hFF;
		16'hFFF1: out_word = 8'hFF;
		16'hFFF2: out_word = 8'hFF;
		16'hFFF3: out_word = 8'hFF;
		16'hFFF4: out_word = 8'hFF;
		16'hFFF5: out_word = 8'hFF;
		16'hFFF6: out_word = 8'hFF;
		16'hFFF7: out_word = 8'hFF;
		16'hFFF8: out_word = 8'h48;
		16'hFFF9: out_word = 8'h45;
		16'hFFFA: out_word = 8'h47;
		16'hFFFB: out_word = 8'h4C;
		16'hFFFC: out_word = 8'h55;
		16'hFFFD: out_word = 8'h4B;
		16'hFFFE: out_word = 8'h56;
		16'hFFFF: out_word = 8'h95;

		default: out_word = 8'hFF;

	endcase

endmodule
