`include "../include/tune.v"

// Pentevo project (c) NedoPC 2010-2011
//
// top module for video output.
//
//
// refactored by TS-Labs

module video_top(

	input  wire        clk, // 28 MHz clock


	// external video outputs
	output wire [ 1:0] vred,
	output wire [ 1:0] vgrn,
	output wire [ 1:0] vblu,
	output wire        vhsync,
	output wire        vvsync,
	output wire        vcsync,


	// aux video inputs
	input  wire [ 5:0] zxborder, // border true color


	// config inputs
	input  wire [ 7:0] vcfg,		// bits 2-0 - vmode:
									//				3'b000 - zx
									//				3'b001 - tiles hi-res
									//				3'b010 - tiles0
									//				3'b011 - tiles0&1
									//				3'b111 - no gfx/border
									// bits 4-3 - raster
									//				2'b0x - 256x192
									//				2'b10 - 320x240
									//				2'b11 - 360x288
									// other bits are described somewhere else


	input  wire        scr_page,   // screen page (bit 3 of 7FFD)

	input  wire        vga_on,     // vga mode ON - scandoubler activated


	// memory synchronization inputs
	input  wire        cbeg,
	input  wire        post_cbeg,
	input  wire        pre_cend,
	input  wire        cend,


	// memory arbiter video port connection
	output wire        video_go,
	output wire [ 1:0] video_bw,
	output wire [20:0] video_addr,
	input  wire [15:0] video_data,
	input  wire        video_strobe,
	input  wire        video_next,

	
	output wire        int_start
);

	// these decoded in video_modedecode.v
	wire mode_zx;
	wire mode_tm;
	wire mode_tp1en;
	wire mode_brd;
	wire mode_pixf_14;
	wire [1:0] rres;


	// synchronization
	wire hsync_start;
	wire line_start;
	wire hint_start;


	wire vblank;
	wire hblank;

	wire vpix;
	wire hpix;

	wire vsync;
	wire hsync;

	wire vga_hsync;

	wire scanin_start;
	wire scanout_start;



	wire fetch_start;
	wire fetch_end;
	wire fetch_sync;


	wire [63:0] pic_bits;


	wire [3:0] pixels;


	wire [5:0] color;
	wire [5:0] vga_color;


	wire [2:0] typos;



	// decode video modes
	video_modedecode video_modedecode(

		.vcfg			(vcfg),

		.mode_zx		(mode_zx),
		.mode_tm		(mode_tm),
		.mode_tp1en		(mode_tp1en),
		.mode_brd		(mode_brd),

		.rres			(rres),

		.mode_pixf_14	(mode_pixf_14),

		.mode_bw		(video_bw)
	);



	// vertical sync generator
	video_sync_v video_sync_v(

		.clk(clk),

		.rres			(rres),

		.hsync_start(hsync_start),
		.line_start(line_start),
		.hint_start(hint_start),

		.vblank(vblank),
		.vsync(vsync),
		.vpix(vpix),
		.vtfetch(vtfetch),

		.int_start(int_start)
	);


	// horizontal sync generator
	video_sync_h video_sync_h(

		.clk(clk),

		.mode_zx		(mode_zx),
		.mode_tm		(mode_tm),
		.mode_brd		(mode_brd),

		.rres			(rres),

		.init			(1'b0),

		.pre_cend		(pre_cend),
		.cend   	 	(cend),


		.hblank			(hblank),
		.hsync			(hsync),
		.hpix			(hpix),

		.line_start		(line_start),
		.hsync_start	(hsync_start),

		.hint_start		(hint_start),

		.scanin_start	(scanin_start),

		.fetch_start	(fetch_start),
		.fetch_end		(fetch_end),
		.tfetch_start	(tfetch_start),
		.tfetch_end		(tfetch_end)

	);


	// address generation
	video_addrgen video_addrgen(

		.clk			(clk),

		.video_addr		(video_addr),
		.video_next		(video_next),

		.line_start		(hsync_start),
		.int_start		(int_start),
		.vpix			(vpix),
		.tfetch			(tfetch),

		.scr_page		(scr_page),

		.mode_zx		(mode_zx),
		.mode_tm		(mode_tm),
		.mode_tp1en		(mode_tp1en),

		);


	// data fetch
	video_fetch video_fetch(

		.clk(clk),

		.pre_cend (pre_cend),
		.cend     (cend    ),

		.vpix(vpix),
		.tfetch			(tfetch),

		.fetch_start(fetch_start),
		.fetch_end  (fetch_end  ),
		.tfetch_start	(tfetch_start),
		.tfetch_end		(tfetch_end),

		.fetch_sync (fetch_sync ),

		.video_data  (video_data  ),
		.video_strobe(video_strobe),
		.video_go    (video_go    ),

		.pic_bits(pic_bits)
	);


	// render fetched data to pixels
	video_render video_render(

		.clk(clk),

		.pic_bits(pic_bits),

		.fetch_sync(fetch_sync),

		.cbeg     (cbeg     ),
		.post_cbeg(post_cbeg),
		.pre_cend (pre_cend ),
		.cend     (cend     ),

		.int_start(int_start),

		.mode_atm_n_pent(mode_atm_n_pent),
		.mode_zx        (mode_zx        ),
		.mode_p_16c     (mode_tm	),
		.mode_p_16c     (mode_tp1en	),
		
		.mode_pixf_14   (mode_pixf_14   ),

		.pixels(pixels)
	);


	// combine border and pixels, apply palette
	video_palframe video_palframe(

		.clk(clk),

		.hblank(hblank),
		.vblank(vblank),

		.hpix(hpix),
		.vpix(vpix),

		.pixels(pixels),
		.border(zxborder),

		.atm_palwr  (atm_palwr  ),
		.atm_paldata(atm_paldata),

		.color(color)
	);


	// VGA hsync doubling
	video_vga_sync_h video_vga_sync_h(

		.clk(clk),

		.hsync_start(hsync_start),

		.scanout_start(scanout_start),

		.vga_hsync(vga_hsync)
	);


	// VGA scandoubling
	video_vga_double video_vga_double(

		.clk(clk),

		.hsync_start  (hsync_start  ),
		.scanout_start(scanout_start),
		.scanin_start (scanin_start ),

		.pix_in(color),

		.pix_out(vga_color)
	);


	// final MUXing of VGA and TV signals
	video_outmux video_outmux(

		.clk(clk),

		.vga_on(vga_on),


		.tvcolor(color),
		.vgacolor(vga_color),

		.vga_hsync(vga_hsync),
		.hsync    (hsync    ),
		.vsync    (vsync    ),

		.vred(vred),
		.vgrn(vgrn),
		.vblu(vblu),

		.vhsync(vhsync),
		.vvsync(vvsync),
		.vcsync(vcsync)
	);






endmodule

