// This module receives 112 MHz as input clock
// and formes strobes for all clocked parts
// (now forms only 28 MHz strobes)

//			0       1       2       3       0       1       2       3       0       1       2       3       
//			0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 
// clk		-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_
// f0		--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__
// q0		--______--______--______--______--______--______--______--______--______--______--______--______
// w0		--______________--______________--______________--______________--______________--______________
// c0		--______________________________--______________________________--______________________________	(ex cbeg)
// c1		________--______________________________--______________________________--______________________	(ex post_cbeg)
// c2		________________--______________________________--______________________________--______________	(ex pre_cend)
// c3		________________________--______________________________--______________________________--______	(ex cend)
// c15		______________________________--______________________________--______________________________--


module clock (

	input wire clk,
	output reg clk175,
	output reg f0, q0, w0, c0, c1, c2, c3, c15

);


	reg [5:0] cnt = 0;

	always @(posedge clk)
		cnt <= cnt + 1;
		
		
	always @*
	begin

		f0 = cnt[0];
		q0 = cnt[1:0] == 2'd0;
		w0 = cnt[2:0] == 3'd0;
		c0 = cnt[3:0] == 4'd0;
		c1 = cnt[3:0] == 4'd4;
		c2 = cnt[3:0] == 4'd8;
		c3 = cnt[3:0] == 4'd12;
		c15 = cnt[3:0] == 4'd15;
		
		clk175 = cnt[5];
		
	end
	

endmodule
