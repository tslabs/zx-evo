`include "../include/tune.v"

// Pentevo project (c) NedoPC 2008-2011
//
// top-level

module top(

	// clocks
	input fclk,
	output clkz_out,
	input clkz_in,

	// z80
	input iorq_n,
	input mreq_n,
	input rd_n,
	input wr_n,
	input m1_n,
	input rfsh_n,
	output int_n,
	output nmi_n,
	output wait_n,
	output res,

	inout [7:0] d,
	input [15:0] a,

	// zxbus and related
	output csrom,
	output romoe_n,
	output romwe_n,

	output rompg0_n,
	output dos_n, // aka rompg1
	output rompg2,
	output rompg3,
	output rompg4,

	input iorqge1,
	input iorqge2,
	output iorq1_n,
	output iorq2_n,

	// DRAM
	inout [15:0] dram_rd,
	output [9:0] dram_ra,
	output rwe_n,
	output rucas_n,
	output rlcas_n,
	output rras0_n,
	output rras1_n,

	// video
	output [1:0] vred,
	output [1:0] vgrn,
	output [1:0] vblu,

	output vhsync,
	output vvsync,
	output vcsync,

	// AY control and audio/tape
	output ay_clk,
	output ay_bdir,
	output ay_bc1,

	output beep,

	// IDE
	output [2:0] ide_a,
	inout [15:0] ide_d,

	output ide_dir,

	input ide_rdy,

	output ide_cs0_n,
	output ide_cs1_n,
	output ide_rs_n,
	output ide_rd_n,
	output ide_wr_n,

	// VG93 and diskdrive
	output vg_clk,

	output vg_cs_n,
	output vg_res_n,

	output vg_hrdy,
	output vg_rclk,
	output vg_rawr,
	output [1:0] vg_a, // disk drive selection
	output vg_wrd,
	output vg_side,

	input step,
	input vg_sl,
	input vg_sr,
	input vg_tr43,
	input rdat_b_n,
	input vg_wf_de,
	input vg_drq,
	input vg_irq,
	input vg_wd,

	// serial links (atmega-fpga, sdcard)
	output sdcs_n,
	output sddo,
	output sdclk,
	input sddi,

	input spics_n,
	input spick,
	input spido,
	output spidi,
	output spiint_n
);

	wire f0, f1, h0, h1, c0, c1, c2, c3;
	wire [1:0] ay_mod;

	clock clock
	(
		.clk(fclk),
		.f0(f0), .f1(f1),
		.h0(h0), .h1(h1),
		.c0(c0), .c1(c1), .c2(c2), .c3(c3),
		.ay_clk(ay_clk),
		.ay_mod(sysconf[4:3])
	);


	wire dos;
	wire vdos;


	wire zpos,zneg;

	wire rst_n; // global reset

	wire [15:0] rddata;

	wire [4:0] rompg = page[4:0];

	wire [7:0] zports_dout;
	wire zports_dataout;
	wire porthit;


	wire [39:0] kbd_data;
	wire [ 7:0] mus_data;
	wire kbd_stb,mus_xstb,mus_ystb,mus_btnstb,kj_stb;

	wire [ 4:0] kbd_port_data;
	wire [ 4:0] kj_port_data;
	wire [ 7:0] mus_port_data;




	wire [7:0] wait_read,wait_write;
	wire wait_rnw;
	wire wait_start_gluclock;
	wire wait_start_comport;
	wire wait_end;
	wire [7:0] gluclock_addr;
	wire [2:0] comport_addr;
	wire [6:0] waits;




	// config signals
	wire [7:0] not_used;
	wire cfg_vga_on;
	wire [1:0] set_nmi;

	// nmi signals
	wire gen_nmi;
	wire clr_nmi;
	wire in_nmi;



	wire tape_in;

	wire [15:0] ideout;
	wire [15:0] idein;
	wire idedataout;


	wire [7:0] zmem_dout;
	wire zmem_dataout;



	wire [7:0] received;
	wire [7:0] tobesent;


	wire intrq,drq;
	wire vg_wrFF;

	wire [1:0] rstrom;




	wire zclk = clkz_in;


	// RESETTER
	wire genrst;

	resetter myrst( .clk(fclk),
	                .rst_in_n(~genrst),
	                .rst_out_n(rst_n) );
	defparam myrst.RST_CNT_SIZE = 6;



	assign nmi_n=gen_nmi ? 1'b0 : 1'bZ;

	assign res= ~rst_n;








	assign ide_rs_n = rst_n;

	assign ide_d = idedataout ? ideout : 16'hZZZZ;
	assign idein = ide_d;

	assign ide_dir = ~idedataout;





	wire [7:0] peff7;


	wire cpm_n;
	wire fnt_wr;



	wire cpu_req,cpu_rnw,cpu_wrbsel,cpu_strobe;
	wire [20:0] cpu_addr;
	// wire [15:0] cpu_rddata;
	wire [7:0] cpu_wrdata;

	wire go;


	wire sd_start;
	wire [7:0] sd_dataout,sd_datain;


	wire tape_read; // data for tapein

	wire beeper_mux; // what is mixed to FPGA beeper output - beeper (0) or tapeout (1)

	wire [2:0] atm_scr_mode;

	wire beeper_wr, covox_wr;


	wire [5:0] palcolor; // palette readback


	wire [1:0] int_turbo;
	wire cpu_next;
	wire cpu_stall;

	wire external_port;


	// fix ATM2-style ROM addressing for PENT-like ROM layout.
	// this causes compications when writing to the flashROM from Z80
	// and need to split and re-build old ATM romfiles before burning in
	// flash
//	wire [1:0] adr_fix;
//	assign adr_fix = ~{ rompg[0], rompg[1] };
//	assign rompg0_n = ~adr_fix[0];
//	assign dos_n    =  adr_fix[1];
//	assign rompg2   =  1'b0;//rompg[2];
//	assign rompg3   =  1'b0;//rompg[3];
//	assign rompg4   =  1'b0;//rompg[4];

	assign rompg0_n = ~rompg[0];
	assign dos_n    =  rompg[1];
	assign rompg2   =  rompg[2];
	assign rompg3   =  rompg[3];
	assign rompg4   =  rompg[4];

	wire zclk_stall;

	zclock zclock
	(
		.fclk(fclk), .rst_n(rst_n), .zclk(zclk), .rfsh_n(rfsh_n), .zclk_out(clkz_out),
		.zpos(zpos), .zneg(zneg),
		.turbo(turbo), .c2(c2), .c0(c0),
		.zclk_stall( cpu_stall | zclk_stall), .int_turbo(int_turbo),
		.external_port(external_port), .iorq_n(iorq_n), .m1_n(m1_n)
	);

    wire [1:0] turbo =  sysconf[1:0];

	wire [7:0] dout_ram;
	wire ena_ram;
	wire [7:0] dout_ports;
	wire ena_ports;


	wire [7:0] border;

	wire drive_ff;


	wire       atm_palwr;
	wire [5:0] atm_paldata;

	wire int_start;


	// data bus out: either RAM data or internal ports data or 0xFF with unused ports
	assign d = ena_ram ? dout_ram : ( ena_ports ? dout_ports : ( drive_ff ? 8'hFF : 8'bZZZZZZZZ ) );




	zbus zxbus( .iorq_n(iorq_n), .rd_n(rd_n), .wr_n(wr_n), .m1_n(m1_n),
	            .iorq1_n(iorq1_n), .iorq2_n(iorq2_n), .iorqge1(iorqge1), .iorqge2(iorqge2),
	            .porthit(porthit), .drive_ff(drive_ff) );



	wire rampage_wr;	    // ports #10AF-#13AF
	wire [7:0] memconf;
	wire [7:0] xt_ramp[0:3];
	wire [7:0] page;
	wire vdos_on, vdos_off;
	wire dos_on, dos_off;
    wire romnram;

    pager pager(
        .clk        (fclk),
        .za         (a),
        .m1         (!m1_n),
        .mreq       (!mreq_n),
        .memconf    (memconf),
        .xt_page    (xt_page),
        .dos        (dos),
        .vdos       (vdos),

        .page       (page),
        .romnram    (romnram),
        .rw_en      (rw_en),
        .dos_on     (dos_on),
        .dos_off    (dos_off),
        .zclk_stall (zclk_stall)

    );



	///////////////////////////
	// DOS signal controller //
	///////////////////////////

	zdos zdos(
	           .fclk(fclk),
			   .rst_n(rst_n),

	           .dos_on  (dos_on),
	           .dos_off (dos_off),
			   .vdos_on (vdos_on),
               .vdos_off(vdos_off),

	           .dos(dos),
	           .vdos(vdos)
	         );




	///////////////////////////
	// Z80 memory controller //
	///////////////////////////

    wire m1_on;
    wire m1_off;

	zmem z80mem
	(
		.fclk (fclk),
		.rst_n(rst_n),

		.zpos(zpos),
		.zneg(zneg),

		.c0    (c0),
		.c1    (c1),
		.c2    (c2),
		.c3    (c3),

		.za    (a),
		.zd_in (d),
		.zd_out(dout_ram),
		.zd_ena(ena_ram),
		.m1_n  (m1_n),
		.rfsh_n(rfsh_n),
		.iorq_n(iorq_n),
		.mreq_n(mreq_n),
		.rd_n  (rd_n),
		.wr_n  (wr_n),

        // .win_page({page[3], page[2], page[1], page[0]}),
		// .win_romnram(romnram),
		.page   (page),
		.romnram(romnram),

		.rw_en(rw_en),
		// .rw_en(1),

		// .rompg  (rompg),
		.romoe_n(romoe_n),
		.romwe_n(romwe_n),
		.csrom  (csrom),

		.vdos_on   (vdos_on),
		.vdos_off  (vdos_off),
        .dos_on    (dos_on),

		.cpu_req   (cpu_req),
		.cpu_rnw   (cpu_rnw),
		.cpu_wrbsel(cpu_wrbsel),
		.cpu_strobe(cpu_strobe),
		.cpu_addr  (cpu_addr),
		.cpu_wrdata(cpu_wrdata),
		// .cpu_rddata(dram_rddata),
		.cpu_rddata(dram_rd),
		.cpu_stall (cpu_stall),
		.cpu_next  (cpu_next),

		.int_turbo(int_turbo)
	);


	wire [20:0] daddr;
	wire dreq;
	wire drnw;
	wire [15:0] dram_rddata;
	wire [15:0] dram_wrdata;
	wire [1:0] dbsel;




	dram dram( .clk(fclk),
	           .rst_n(rst_n),

	           .addr(daddr),
	           .req(dreq),
	           .rnw(drnw),
	           .c0(c0),
	           .c1(c1),
	           .c2(c2),
	           .c3(c3),
	           .rddata(dram_rddata),
	           .wrdata(dram_wrdata),
	           .bsel(dbsel),

	           .ra(dram_ra),
	           .rd(dram_rd),
	           .rwe_n(rwe_n),
	           .rucas_n(rucas_n),
	           .rlcas_n(rlcas_n),
	           .rras0_n(rras0_n),
	           .rras1_n(rras1_n)
	         );


	wire [4:0] video_bw;

	wire [20:0] video_addr;
	wire video_strobe;
	wire video_next;

	wire [20:0] dma_addr;
	wire [15:0] dma_wrdata;
	wire dma_req;
	wire dma_rnw;
	wire dma_next;
	wire dma_strobe;

	wire [20:0] ts_addr;
	wire ts_req;
	wire ts_next;

	arbiter dramarb(
					 .clk(fclk),
	                 .c2(c2),
	                 .c3(c3),

	                 .rst_n(rst_n),

	                 .dram_addr(daddr),
	                 .dram_req(dreq),
	                 .dram_rnw(drnw),
	                 .dram_bsel(dbsel),
	                 .dram_wrdata(dram_wrdata),

	                 //.cpu_waitcyc(cpu_waitcyc),
	                 .cpu_addr		(cpu_addr),
	                 .cpu_wrdata	(cpu_wrdata),
	                 .cpu_req		(cpu_req),
	                 .cpu_rnw		(cpu_rnw),
	                 .cpu_wrbsel	(cpu_wrbsel),
					 .cpu_next		(cpu_next),
	                 .cpu_strobe	(cpu_strobe),

	                 .go(go),
	                 .video_bw(video_bw),
	                 .video_addr(video_addr),
	                 .video_strobe(video_strobe),
	                 .video_next(video_next),

	                 .dma_addr		(dma_addr),
	                 .dma_wrdata	(dma_wrdata),
	                 .dma_req		(dma_req),
	                 .dma_rnw		(dma_rnw),
					 .dma_next		(dma_next),

					 .ts_req		(ts_req),
					 .ts_addr		(ts_addr),
					 .ts_next		(ts_next)
	);


        wire border_wr   ;
        wire zborder_wr  ;
        wire zvpage_wr	 ;
        wire vpage_wr	 ;
        wire vconf_wr	 ;
        wire x_offsl_wr	 ;
        wire x_offsh_wr	 ;
        wire y_offsl_wr	 ;
        wire y_offsh_wr	 ;
        wire palsel_wr	 ;
        wire hint_beg_wr ;
        wire vint_begl_wr;
        wire vint_begh_wr;
        wire tsconf_wr	 ;
        wire tmpage_wr	 ;
        wire t0gpage_wr	 ;
        wire t1gpage_wr	 ;
        wire sgpage_wr	 ;

    // wire [1:0] vred0;
    // assign vred = vred0 | {2{t}};

	video_top video_top(

		.clk(fclk),
		.zclk(zclk),
        .res(res),
		.f0(f0), .f1(f1),
		.h0(h0), .h1(h1),
		.c0(c0), .c1(c1), .c2(c2), .c3(c3),
		// .t(t),	//debug!!!

		.vred(vred),
		.vgrn(vgrn),
		.vblu(vblu),
		.hsync(vhsync),
		.vsync(vvsync),
		.csync(vcsync),

		.vga_on(cfg_vga_on),

        .border_wr      (border_wr),
        .zborder_wr     (zborder_wr),
		.zvpage_wr	    (zvpage_wr),
		.vpage_wr	    (vpage_wr),
		.vconf_wr	    (vconf_wr),
		.x_offsl_wr	    (x_offsl_wr),
		.x_offsh_wr	    (x_offsh_wr),
		.y_offsl_wr	    (y_offsl_wr),
		.y_offsh_wr	    (y_offsh_wr),
		.palsel_wr	    (palsel_wr),
		.hint_beg_wr    (hint_beg_wr),
		.vint_begl_wr   (vint_begl_wr),
		.vint_begh_wr   (vint_begh_wr),
		.tsconf_wr	    (tsconf_wr),
		.tmpage_wr	    (tmpage_wr),
		.t0gpage_wr	    (t0gpage_wr),
		.t1gpage_wr	    (t1gpage_wr),
		.sgpage_wr	    (sgpage_wr),

		.video_addr     (video_addr),
		.video_bw		(video_bw),
		.video_go       (go),
		.dram_rddata    (dram_rddata),      // reg'ed, should be latched by c3
   		.dram_rdata     (dram_rd),               // raw, should be latched by c2
		.video_strobe   (video_strobe),
		.video_next     (video_next),

		.ts_req			(ts_req),
		.ts_addr		(ts_addr),
		.ts_next		(ts_next),

		.a(a), .d(d),
		.cram_data_in({d[6:0], zmd}),
		.sfys_data_in({d[7:0], zmd}),
		.cram_we(cram_we),
		.sfys_we(sfys_we),
		.int_start(int_start)

	);


	slavespi slavespi(
		.fclk(fclk), .rst_n(rst_n),

		.spics_n(spics_n), .spidi(spidi),
		.spido(spido), .spick(spick),
		.status_in({/* wait_rnw */ wr_n, waits[6:0]}), .genrst(genrst),
		.rstrom(rstrom), .kbd_out(kbd_data),
		.kbd_stb(kbd_stb), .mus_out(mus_data),
		.mus_xstb(mus_xstb), .mus_ystb(mus_ystb),
		.mus_btnstb(mus_btnstb), .kj_stb(kj_stb),
		.gluclock_addr(gluclock_addr),
		.comport_addr (comport_addr),
		.wait_write(wait_write),
		.wait_read(wait_read),
		.wait_rnw(wait_rnw),
		.wait_end(wait_end),
		.config0( { not_used[7:4], beeper_mux, tape_read, set_nmi[0], cfg_vga_on} )
	);

	zkbdmus zkbdmus( .fclk(fclk), .rst_n(rst_n),
	                 .kbd_in(kbd_data), .kbd_stb(kbd_stb),
	                 .mus_in(mus_data), .mus_xstb(mus_xstb),
	                 .mus_ystb(mus_ystb), .mus_btnstb(mus_btnstb),
	                 .kj_stb(kj_stb), .kj_data(kj_port_data),
	                 .zah(a[15:8]), .kbd_data(kbd_port_data),
	                 .mus_data(mus_port_data)
	               );


		wire [7:0]	   zmd	;

    zmaps zmaps(
				.zclk   (zclk),
				.mreq_n (mreq_n),
				.wr_n   (wr_n),
				.a      (a),
				.d      (d),
				.fmaddr (fmaddr),
				.zmd    (zmd),
				.cram_we(cram_we),
				.sfys_we(sfys_we)
				);


	wire rst;
	wire iorq;
	wire iorq_s;
	wire mreq;
	wire m1;
	wire rd;
	wire wr;
	wire rdwr;
	wire iord;
	wire iowr;
	wire iorw;
	wire memrd;
	wire memwr;
	wire memrw;

    zsignals zsignals(
                .clk    (fclk),
				.zclk   (zclk),

				.rst_n  (rst_n),

                .iorq_n (iorq_n),
                .mreq_n (mreq_n),
                .m1_n   (m1_n),
                .rd_n   (rd_n),
                .wr_n   (wr_n),

                .rst    (rst),
                .iorq   (iorq),
                .iorq_s (iorq_s),
                .mreq   (mreq),
                .m1     (m1),
                .rd     (rd),
                .wr     (wr),
                .rdwr   (rdwr),
                .iord   (iord),
                .iowr   (iowr),
                .iorw   (iorw),
                .memrd  (memrd),
                .memwr  (memwr),
                .memrw  (memrw)
                );


		wire cram_we;
		wire sfys_we;


		wire [31:0] xt_page;

		wire [8:0] dmaport_wr;
		wire [4:0] fmaddr;

		wire [7:0] sysconf;
		wire [7:0] im2vect ;
		wire [3:0] fddvirt ;

	zports zports(
                    .zclk(zclk), .fclk(fclk),
                    .zpos(zpos), .zneg(zneg),
                    .din(d), .dout(dout_ports), .dataout(ena_ports),
                    .a(a),

                    .rst_n(rst_n),
                    .iorq_n(iorq_n),
                    .mreq_n(mreq_n),
                    .m1_n(m1_n),
                    .rd_n(rd_n),
                    .wr_n(wr_n),

                    .iorq(iorq),
                    .iorq_s(iorq_s),
                    .mreq(mreq),
                    .m1(m1),
                    .iord(iord),
                    .iowr(iowr),
                    .iorw(iorw),
                    .rd(rd),
                    .wr(wr),
                    .rdwr(rdwr),

                    .porthit(porthit),
                    .ay_bdir(ay_bdir), .ay_bc1(ay_bc1),
                    .peff7(peff7),
                    .rstrom(rstrom), .vg_intrq(intrq), .vg_drq(drq), .vg_wrFF(vg_wrFF), .vg_cs_n(vg_cs_n),
                    .sd_start(sd_start), .sd_dataout(sd_dataout), .sd_datain(sd_datain), .sdcs_n(sdcs_n),
                    .idein(idein), .ideout(ideout), .idedataout(idedataout),
                    .ide_a(ide_a), .ide_cs0_n(ide_cs0_n), .ide_cs1_n(ide_cs1_n),
                    .ide_wr_n(ide_wr_n), .ide_rd_n(ide_rd_n),

                    .border_wr      (border_wr),
                    .zborder_wr     (zborder_wr),
					.zvpage_wr	    (zvpage_wr),
					.vpage_wr	    (vpage_wr),
					.vconf_wr	    (vconf_wr),
					.x_offsl_wr	    (x_offsl_wr),
					.x_offsh_wr	    (x_offsh_wr),
					.y_offsl_wr	    (y_offsl_wr),
					.y_offsh_wr	    (y_offsh_wr),
					.palsel_wr	    (palsel_wr),
					.hint_beg_wr    (hint_beg_wr),
					.vint_begl_wr   (vint_begl_wr),
					.vint_begh_wr   (vint_begh_wr),
					.tsconf_wr	    (tsconf_wr),
					.tmpage_wr	    (tmpage_wr),
					.t0gpage_wr	    (t0gpage_wr),
					.t1gpage_wr	    (t1gpage_wr),
					.sgpage_wr	    (sgpage_wr),

					.xt_page (xt_page),

					.fmaddr		(fmaddr),

					.sysconf	(sysconf),
					.memconf	(memconf),
					.im2vect	(im2vect),
					.fddvirt	(fddvirt),
                    .vg_a       (vg_a),
                    .dos        (dos),
                    .vdos       (vdos),
                    .vdos_on    (vdos_on),
                    .vdos_off   (vdos_off),

					.dmaport_wr (dmaport_wr),
                    .dma_act	(dma_act),

                    .keys_in(kbd_port_data),
                    .mus_in (mus_port_data),
                    .kj_in  (kj_port_data),

                    .tape_read(tape_read),

                    .gluclock_addr(gluclock_addr),
                    .comport_addr (comport_addr),
                    .wait_start_gluclock(wait_start_gluclock),
                    .wait_start_comport (wait_start_comport),
                    .wait_rnw  (wait_rnw),
                    .wait_write(wait_write),
`ifndef SIMULATE
                    .wait_read (wait_read),
`else
                    .wait_read(8'hFF),
`endif
					.beeper_wr(beeper_wr),
					.covox_wr (covox_wr),

					.fnt_wr(fnt_wr),
					.clr_nmi(clr_nmi),


					// .pages(~{ rd_pages[7], rd_pages[6],
							// rd_pages[5], rd_pages[4],
							// rd_pages[3], rd_pages[2],
							// rd_pages[1], rd_pages[0] }),

					// .ramnroms( rd_ramnrom),
					// .dos7ffds( rd_dos7ffd),

					.external_port(external_port)

					// .set_nmi(set_nmi[1])
	);


	wire dma_act;
	wire dma_wait;

	dma dma(
		.clk		(fclk),
		.c2		    (c2),
        .rst_n		(rst_n),

		.zdata		(d),
		.dmaport_wr	(dmaport_wr),
		.dma_act	(dma_act),
		.dma_wait	(dma_wait),
		.rfsh_n     (rfsh_n),

		.dram_addr	(dma_addr),
		.dram_rnw	(dma_rnw),
		.dram_req	(dma_req),
		.dram_rddata(dram_rd),
		.dram_wrdata(dma_wrdata),
		.dram_next	(dma_next)
	);


	zint zint(
		.fclk(fclk),
		.zpos(zpos),
		.zneg(zneg),

		.int_start(int_start),
		.vdos(vdos),

		.iorq_n(iorq_n),
		.m1_n  (m1_n),

		.int_n(int_n)
	);

	znmi znmi(
		.rst_n(rst_n),
		.fclk(fclk),
		.zpos(zpos),
		.zneg(zneg),

		.rfsh_n(rfsh_n),

		.int_start(int_start),

		.set_nmi(set_nmi),
		.clr_nmi(clr_nmi),

		.in_nmi (in_nmi),
		.gen_nmi(gen_nmi)
	);




	zwait zwait(
                 .wait_start_gluclock(wait_start_gluclock),
	             .wait_start_comport (wait_start_comport),
	             .wait_end(wait_end),
	             .rst_n(rst_n),
                 .dma_wait(dma_wait),
	             .wait_n(wait_n),
	             .waits(waits),
	             .spiint_n(spiint_n)
    );




	// wire [1:0] vg_ddrv;
	// assign vg_a[0] = vg_ddrv[0] ? 1'b1 : 1'b0; // possibly open drain?
	// assign vg_a[1] = vg_ddrv[1] ? 1'b1 : 1'b0;

	vg93 vgshka( .zclk(zclk), .rst_n(rst_n), .fclk(fclk), .vg_clk(vg_clk),
	             .vg_res_n(vg_res_n), .din(d), .intrq(intrq), .drq(drq), .vg_wrFF(vg_wrFF),
	             .vg_hrdy(vg_hrdy), .vg_rclk(vg_rclk), .vg_rawr(vg_rawr),
	             .vg_wrd(vg_wrd), .vg_side(vg_side), .step(step), .vg_sl(vg_sl), .vg_sr(vg_sr),
	             .vg_tr43(vg_tr43), .rdat_n(rdat_b_n), .vg_wf_de(vg_wf_de), .vg_drq(vg_drq),
	             .vg_irq(vg_irq), .vg_wd(vg_wd) );




	spi2 zspi( .clk(fclk), .sck(sdclk), .sdo(sddo), .sdi(sddi), .start(sd_start),
	           .speed(2'b00),	// this is 14 MHz at 28 Mhz Altera clock
			   .din(sd_datain), .dout(sd_dataout) );





	  //////////////////////////////////////
	 // sound: beeper, tapeout and covox //
	//////////////////////////////////////

	sound sound(

		.clk(fclk), .f0(f0),

		.din(d),

		.beeper_wr(beeper_wr),
		.covox_wr (covox_wr),

		.beeper_mux(beeper_mux),

		.sound_bit(beep)
	);


endmodule

