
`include "../include/tune.v"

module rom(
	input wire [15:0] a,
	output reg [7:0] d

);


	always @*
	case (a)
16'h0000:	d = 8'hF3;	// di
16'h0001:	d = 8'h01;  // ld bc, #FE
16'h0002:	d = 8'hFE;  //
16'h0003:	d = 8'h00;  //
16'h0004:	d = 8'h3C;	// inc a
16'h0005:	d = 8'hED;	// out (c), a
16'h0006:	d = 8'h79;	//
16'h0007:	d = 8'h18;  // jr #0004
16'h0008:	d = 8'hFB;	//
16'h0009:	d = 8'h00;	//
16'h000A:	d = 8'h00;	//
16'h000B:	d = 8'h00;	//
16'h000C:	d = 8'h00;	//
16'h000D:	d = 8'h00;	//
16'h000E:	d = 8'h00;	//
16'h000F:	d = 8'h00;	//
16'h0010:	d = 8'h04;	// rubbish
16'h0011:	d = 8'h15;	//
16'h0012:	d = 8'h63;	//
16'h0013:	d = 8'hD5;	//
16'h0014:	d = 8'h12;	//
16'h0015:	d = 8'hF7;	//
16'h0016:	d = 8'h91;	//
16'h0017:	d = 8'hD9;	//
16'h0018:	d = 8'hA9;	//
16'h0019:	d = 8'h12;	//
16'h001A:	d = 8'hA8;	//
16'h001B:	d = 8'h46;	//
16'h001C:	d = 8'h66;	//
16'h001D:	d = 8'h0D;	//
16'h001E:	d = 8'hA5;	//
16'h001F:	d = 8'h13;	//
16'h0020:	d = 8'hA9;	//
16'h0021:	d = 8'h5E;	//
16'h0022:	d = 8'hD2;	//
16'h0023:	d = 8'h2C;	//
16'h0024:	d = 8'hAD;	//
16'h0025:	d = 8'h79;	//
16'h0026:	d = 8'h74;	//
16'h0027:	d = 8'h36;	//
16'h0028:	d = 8'h3F;	//
16'h0029:	d = 8'h3A;	//
16'h002A:	d = 8'h5D;	//
16'h002B:	d = 8'h59;	//
16'h002C:	d = 8'h9E;	//
16'h002D:	d = 8'hAA;	//
16'h002E:	d = 8'hC8;	//
16'h002F:	d = 8'hFF;	//
16'h0030:	d = 8'hD3;	//
16'h0031:	d = 8'h5A;	//
16'h0032:	d = 8'hFE;	//
16'h0033:	d = 8'h79;	//
16'h0034:	d = 8'h4B;	//
16'h0035:	d = 8'hD9;	//
16'h0036:	d = 8'h8F;	//
16'h0037:	d = 8'h55;	//
16'h0038:	d = 8'hCF;	//
16'h0039:	d = 8'h53;	//
16'h003A:	d = 8'h5C;	//
16'h003B:	d = 8'hAD;	//
16'h003C:	d = 8'h0A;	//
16'h003D:	d = 8'h22;	//
16'h003E:	d = 8'h7B;	//
16'h003F:	d = 8'h18;	//
16'h0040:	d = 8'h12;	//
16'h0041:	d = 8'h87;	//
16'h0042:	d = 8'h09;	//
16'h0043:	d = 8'hD1;	//
16'h0044:	d = 8'hB8;	//
16'h0045:	d = 8'hA0;	//
16'h0046:	d = 8'h57;	//
16'h0047:	d = 8'h50;	//
16'h0048:	d = 8'hC7;	//
16'h0049:	d = 8'h82;	//
16'h004A:	d = 8'h12;	//
16'h004B:	d = 8'hAE;	//
16'h004C:	d = 8'hB0;	//
16'h004D:	d = 8'h6D;	//
16'h004E:	d = 8'h30;	//
16'h004F:	d = 8'hB2;	//
16'h0050:	d = 8'h2B;	//
16'h0051:	d = 8'hCA;	//
16'h0052:	d = 8'h54;	//
16'h0053:	d = 8'h8F;	//
16'h0054:	d = 8'hCF;	//
16'h0055:	d = 8'hB5;	//
16'h0056:	d = 8'h38;	//
16'h0057:	d = 8'hF2;	//
16'h0058:	d = 8'hF8;	//
16'h0059:	d = 8'h2A;	//
16'h005A:	d = 8'hE2;	//
16'h005B:	d = 8'h00;	//
16'h005C:	d = 8'h25;	//
16'h005D:	d = 8'h01;	//
16'h005E:	d = 8'hC5;	//
16'h005F:	d = 8'hC4;	//
16'h0060:	d = 8'h90;	//
16'h0061:	d = 8'h55;	//
16'h0062:	d = 8'h8A;	//
16'h0063:	d = 8'h2C;	//
16'h0064:	d = 8'h60;	//
16'h0065:	d = 8'h50;	//
16'h0066:	d = 8'h34;	//
16'h0067:	d = 8'h91;	//
16'h0068:	d = 8'h09;	//
16'h0069:	d = 8'h29;	//
16'h006A:	d = 8'h40;	//
16'h006B:	d = 8'h58;	//
16'h006C:	d = 8'h9C;	//
16'h006D:	d = 8'hF1;	//
16'h006E:	d = 8'h08;	//
16'h006F:	d = 8'h4A;	//
16'h0070:	d = 8'h26;	//
16'h0071:	d = 8'h54;	//
16'h0072:	d = 8'h27;	//
16'h0073:	d = 8'h15;	//
16'h0074:	d = 8'h97;	//
16'h0075:	d = 8'h58;	//
16'h0076:	d = 8'hE9;	//
16'h0077:	d = 8'h2A;	//
16'h0078:	d = 8'h33;	//
16'h0079:	d = 8'h24;	//
16'h007A:	d = 8'h42;	//
16'h007B:	d = 8'hBA;	//
16'h007C:	d = 8'h64;	//
16'h007D:	d = 8'hC3;	//
16'h007E:	d = 8'h64;	//
16'h007F:	d = 8'hE4;	//
16'h0080:	d = 8'hE9;	//
16'h0081:	d = 8'h48;	//
16'h0082:	d = 8'hE3;	//
16'h0083:	d = 8'h6F;	//
16'h0084:	d = 8'h44;	//
16'h0085:	d = 8'h05;	//
16'h0086:	d = 8'h26;	//
16'h0087:	d = 8'h4B;	//
16'h0088:	d = 8'h3F;	//
16'h0089:	d = 8'h66;	//
16'h008A:	d = 8'h0C;	//
16'h008B:	d = 8'hEC;	//
16'h008C:	d = 8'hE0;	//
16'h008D:	d = 8'h70;	//
16'h008E:	d = 8'h95;	//
16'h008F:	d = 8'hFF;	//
16'h0090:	d = 8'hF3;	//
16'h0091:	d = 8'h70;	//
16'h0092:	d = 8'h64;	//
16'h0093:	d = 8'hFD;	//
16'h0094:	d = 8'h15;	//
16'h0095:	d = 8'h0D;	//
16'h0096:	d = 8'h89;	//
16'h0097:	d = 8'h1A;	//
16'h0098:	d = 8'h12;	//
16'h0099:	d = 8'h6B;	//
16'h009A:	d = 8'h09;	//
16'h009B:	d = 8'h16;	//
16'h009C:	d = 8'h03;	//
16'h009D:	d = 8'h48;	//
16'h009E:	d = 8'h4E;	//
16'h009F:	d = 8'hDB;	//
16'h00A0:	d = 8'h8A;	//
16'h00A1:	d = 8'h1D;	//
16'h00A2:	d = 8'h2A;	//
16'h00A3:	d = 8'h80;	//
16'h00A4:	d = 8'hD9;	//
16'h00A5:	d = 8'h42;	//
16'h00A6:	d = 8'h98;	//
16'h00A7:	d = 8'hAB;	//
16'h00A8:	d = 8'h38;	//
16'h00A9:	d = 8'h46;	//
16'h00AA:	d = 8'h4E;	//
16'h00AB:	d = 8'h4C;	//
16'h00AC:	d = 8'h88;	//
16'h00AD:	d = 8'hEA;	//
16'h00AE:	d = 8'h1D;	//
16'h00AF:	d = 8'h42;	//
16'h00B0:	d = 8'h59;	//
16'h00B1:	d = 8'hA8;	//
16'h00B2:	d = 8'h86;	//
16'h00B3:	d = 8'h8C;	//
16'h00B4:	d = 8'hB0;	//
16'h00B5:	d = 8'h80;	//
16'h00B6:	d = 8'h96;	//
16'h00B7:	d = 8'h32;	//
16'h00B8:	d = 8'h2B;	//
16'h00B9:	d = 8'h4D;	//
16'h00BA:	d = 8'h35;	//
16'h00BB:	d = 8'h08;	//
16'h00BC:	d = 8'h6E;	//
16'h00BD:	d = 8'hD9;	//
16'h00BE:	d = 8'h14;	//
16'h00BF:	d = 8'h25;	//
16'h00C0:	d = 8'h0C;	//
16'h00C1:	d = 8'hA5;	//
16'h00C2:	d = 8'h69;	//
16'h00C3:	d = 8'h63;	//
16'h00C4:	d = 8'h59;	//
16'h00C5:	d = 8'h2D;	//
16'h00C6:	d = 8'h30;	//
16'h00C7:	d = 8'h56;	//
16'h00C8:	d = 8'h7C;	//
16'h00C9:	d = 8'hCA;	//
16'h00CA:	d = 8'h46;	//
16'h00CB:	d = 8'h95;	//
16'h00CC:	d = 8'h46;	//
16'h00CD:	d = 8'hB3;	//
16'h00CE:	d = 8'h27;	//
16'h00CF:	d = 8'h22;	//
16'h00D0:	d = 8'hDC;	//
16'h00D1:	d = 8'h0B;	//
16'h00D2:	d = 8'h51;	//
16'h00D3:	d = 8'h48;	//
16'h00D4:	d = 8'h41;	//
16'h00D5:	d = 8'h94;	//
16'h00D6:	d = 8'h2E;	//
16'h00D7:	d = 8'hA3;	//
16'h00D8:	d = 8'h2A;	//
16'h00D9:	d = 8'hDD;	//
16'h00DA:	d = 8'hB9;	//
16'h00DB:	d = 8'h84;	//
16'h00DC:	d = 8'h43;	//
16'h00DD:	d = 8'hE6;	//
16'h00DE:	d = 8'h84;	//
16'h00DF:	d = 8'h82;	//
16'h00E0:	d = 8'hB8;	//
16'h00E1:	d = 8'h7D;	//
16'h00E2:	d = 8'hBF;	//
16'h00E3:	d = 8'hC8;	//
16'h00E4:	d = 8'hD7;	//
16'h00E5:	d = 8'h9C;	//
16'h00E6:	d = 8'hFF;	//
16'h00E7:	d = 8'h4C;	//
16'h00E8:	d = 8'h53;	//
16'h00E9:	d = 8'h80;	//
16'h00EA:	d = 8'h0E;	//
16'h00EB:	d = 8'hD6;	//
16'h00EC:	d = 8'h15;	//
16'h00ED:	d = 8'h22;	//
16'h00EE:	d = 8'h8B;	//
16'h00EF:	d = 8'h88;	//
16'h00F0:	d = 8'h4D;	//
16'h00F1:	d = 8'h19;	//
16'h00F2:	d = 8'hC2;	//
16'h00F3:	d = 8'hC0;	//
16'h00F4:	d = 8'hCC;	//
16'h00F5:	d = 8'hE6;	//
16'h00F6:	d = 8'h70;	//
16'h00F7:	d = 8'h21;	//
16'h00F8:	d = 8'h44;	//
16'h00F9:	d = 8'h32;	//
16'h00FA:	d = 8'h02;	//
16'h00FB:	d = 8'h49;	//
16'h00FC:	d = 8'hF2;	//
16'h00FD:	d = 8'hBD;	//
16'h00FE:	d = 8'h17;	//
16'h00FF:	d = 8'h32;	//
16'h0100:	d = 8'hAB;	//
16'h0101:	d = 8'hBF;  //
16'h0102:	d = 8'h61;  //
16'h0103:	d = 8'h80;  //
16'h0104:	d = 8'hEC;	//
16'h0105:	d = 8'hBD;	//
16'h0106:	d = 8'hA3;	//
16'h0107:	d = 8'hD1;  //
16'h0108:	d = 8'hE4;	//
16'h0109:	d = 8'h53;	//
16'h010A:	d = 8'h11;	//
16'h010B:	d = 8'h08;	//
16'h010C:	d = 8'hCA;	//
16'h010D:	d = 8'h4B;	//
16'h010E:	d = 8'h02;	//
16'h010F:	d = 8'h49;	//
16'h0110:	d = 8'hEF;	//
16'h0111:	d = 8'h13;	//
16'h0112:	d = 8'h44;	//
16'h0113:	d = 8'h95;	//
16'h0114:	d = 8'h97;	//
16'h0115:	d = 8'hC5;	//
16'h0116:	d = 8'h64;	//
16'h0117:	d = 8'h25;	//
16'h0118:	d = 8'h09;	//
16'h0119:	d = 8'hDE;	//
16'h011A:	d = 8'h4E;	//
16'h011B:	d = 8'h59;	//
16'h011C:	d = 8'h19;	//
16'h011D:	d = 8'hD2;	//
16'h011E:	d = 8'h26;	//
16'h011F:	d = 8'h84;	//
16'h0120:	d = 8'h64;	//
16'h0121:	d = 8'h6D;	//
16'h0122:	d = 8'h2A;	//
16'h0123:	d = 8'h88;	//
16'h0124:	d = 8'h51;	//
16'h0125:	d = 8'h08;	//
16'h0126:	d = 8'h8F;	//
16'h0127:	d = 8'hEA;	//
16'h0128:	d = 8'h1B;	//
16'h0129:	d = 8'h40;	//
16'h012A:	d = 8'h81;	//
16'h012B:	d = 8'h34;	//
16'h012C:	d = 8'h3D;	//
16'h012D:	d = 8'h64;	//
16'h012E:	d = 8'h96;	//
16'h012F:	d = 8'h28;	//
16'h0130:	d = 8'h60;	//
16'h0131:	d = 8'h52;	//
16'h0132:	d = 8'h61;	//
16'h0133:	d = 8'hA1;	//
16'h0134:	d = 8'hC4;	//
16'h0135:	d = 8'h10;	//
16'h0136:	d = 8'h68;	//
16'h0137:	d = 8'h50;	//
16'h0138:	d = 8'h05;	//
16'h0139:	d = 8'h30;	//
16'h013A:	d = 8'h7D;	//
16'h013B:	d = 8'hFF;	//
16'h013C:	d = 8'hF3;	//
16'h013D:	d = 8'h72;	//
16'h013E:	d = 8'h64;	//
16'h013F:	d = 8'hF5;	//
16'h0140:	d = 8'h14;	//
16'h0141:	d = 8'hCD;	//
16'h0142:	d = 8'h7D;	//
16'h0143:	d = 8'h1A;	//
16'h0144:	d = 8'h01;	//
16'h0145:	d = 8'h69;	//
16'h0146:	d = 8'h89;	//
16'h0147:	d = 8'h40;	//
16'h0148:	d = 8'h80;	//
16'h0149:	d = 8'h00;	//
16'h014A:	d = 8'h03;	//
16'h014B:	d = 8'h48;	//
16'h014C:	d = 8'h02;	//
16'h014D:	d = 8'hA4;	//
16'h014E:	d = 8'h5C;	//
16'h014F:	d = 8'h84;	//
16'h0150:	d = 8'h13;	//
16'h0151:	d = 8'h43;	//
16'h0152:	d = 8'h4E;	//
16'h0153:	d = 8'h9A;	//
16'h0154:	d = 8'h4C;	//
16'h0155:	d = 8'h0B;	//
16'h0156:	d = 8'h93;	//
16'h0157:	d = 8'h2E;	//
16'h0158:	d = 8'h33;	//
16'h0159:	d = 8'hAF;	//
16'h015A:	d = 8'h24;	//
16'h015B:	d = 8'hA8;	//
16'h015C:	d = 8'h3C;	//
16'h015D:	d = 8'hF9;	//
16'h015E:	d = 8'h7C;	//
16'h015F:	d = 8'h6D;	//
16'h0160:	d = 8'h04;	//
16'h0161:	d = 8'h57;	//
16'h0162:	d = 8'h59;	//
16'h0163:	d = 8'h35;	//
16'h0164:	d = 8'h5B;	//
16'h0165:	d = 8'h83;	//
16'h0166:	d = 8'h05;	//
16'h0167:	d = 8'h55;	//
16'h0168:	d = 8'h72;	//
16'h0169:	d = 8'h15;	//
16'h016A:	d = 8'hDC;	//
16'h016B:	d = 8'hA4;	//
16'h016C:	d = 8'hCA;	//
16'h016D:	d = 8'hBA;	//
16'h016E:	d = 8'hED;	//
16'h016F:	d = 8'h64;	//
16'h0170:	d = 8'h48;	//
16'h0171:	d = 8'h8A;	//
16'h0172:	d = 8'hD0;	//
16'h0173:	d = 8'hD1;	//
16'h0174:	d = 8'h02;	//
16'h0175:	d = 8'h06;	//
16'h0176:	d = 8'h4F;	//
16'h0177:	d = 8'h91;	//
16'h0178:	d = 8'h1C;	//
16'h0179:	d = 8'h40;	//
16'h017A:	d = 8'h92;	//
16'h017B:	d = 8'hBB;	//
16'h017C:	d = 8'h44;	//
16'h017D:	d = 8'h0D;	//
16'h017E:	d = 8'hA0;	//
16'h017F:	d = 8'h24;	//
16'h0180:	d = 8'h39;	//
16'h0181:	d = 8'hE9;	//
16'h0182:	d = 8'hB2;	//
16'h0183:	d = 8'h45;	//
16'h0184:	d = 8'hB2;	//
16'h0185:	d = 8'h97;	//
16'h0186:	d = 8'h5F;	//
16'h0187:	d = 8'hBA;	//
16'h0188:	d = 8'hBD;	//
16'h0189:	d = 8'h36;	//
16'h018A:	d = 8'h7D;	//
16'h018B:	d = 8'hB9;	//
16'h018C:	d = 8'hFA;	//
16'h018D:	d = 8'hB8;	//
16'h018E:	d = 8'h13;	//
16'h018F:	d = 8'hC0;	//
16'h0190:	d = 8'hFB;	//
16'h0191:	d = 8'hCB;	//
16'h0192:	d = 8'h22;	//
16'h0193:	d = 8'hB2;	//
16'h0194:	d = 8'h5F;	//
16'h0195:	d = 8'hD0;	//
16'h0196:	d = 8'hB7;	//
16'h0197:	d = 8'hA9;	//
16'h0198:	d = 8'hEF;	//
16'h0199:	d = 8'h60;	//
16'h019A:	d = 8'h91;	//
16'h019B:	d = 8'h5E;	//
16'h019C:	d = 8'hF2;	//
16'h019D:	d = 8'hE9;	//
16'h019E:	d = 8'hE7;	//
16'h019F:	d = 8'h9E;	//
16'h01A0:	d = 8'hD1;	//
16'h01A1:	d = 8'hED;	//
16'h01A2:	d = 8'h61;	//
16'h01A3:	d = 8'h50;	//
16'h01A4:	d = 8'h4A;	//
16'h01A5:	d = 8'h09;	//
16'h01A6:	d = 8'h9C;	//
16'h01A7:	d = 8'hE0;	//
16'h01A8:	d = 8'h31;	//
16'h01A9:	d = 8'hC4;	//
16'h01AA:	d = 8'h17;	//
16'h01AB:	d = 8'h0A;	//
16'h01AC:	d = 8'hCA;	//
16'h01AD:	d = 8'h85;	//
16'h01AE:	d = 8'hC4;	//
16'h01AF:	d = 8'h50;	//
16'h01B0:	d = 8'h97;	//
16'h01B1:	d = 8'h80;	//
16'h01B2:	d = 8'hB4;	//
16'h01B3:	d = 8'h08;	//
16'h01B4:	d = 8'hD2;	//
16'h01B5:	d = 8'h9C;	//
16'h01B6:	d = 8'hB4;	//
16'h01B7:	d = 8'h6D;	//
16'h01B8:	d = 8'hDA;	//
16'h01B9:	d = 8'h50;	//
16'h01BA:	d = 8'hDD;	//
16'h01BB:	d = 8'hE9;	//
16'h01BC:	d = 8'h6B;	//
16'h01BD:	d = 8'hBD;	//
16'h01BE:	d = 8'h30;	//
16'h01BF:	d = 8'hC4;	//
16'h01C0:	d = 8'h3F;	//
16'h01C1:	d = 8'h2E;	//
16'h01C2:	d = 8'hAB;	//
16'h01C3:	d = 8'h4F;	//
16'h01C4:	d = 8'h62;	//
16'h01C5:	d = 8'hE5;	//
16'h01C6:	d = 8'h4A;	//
16'h01C7:	d = 8'hB0;	//
16'h01C8:	d = 8'h28;	//
16'h01C9:	d = 8'hE2;	//
16'h01CA:	d = 8'hD1;	//
16'h01CB:	d = 8'h8A;	//
16'h01CC:	d = 8'h9D;	//
16'h01CD:	d = 8'hE3;	//
16'h01CE:	d = 8'h4D;	//
16'h01CF:	d = 8'hC3;	//
16'h01D0:	d = 8'h4C;	//
16'h01D1:	d = 8'h0E;	//
16'h01D2:	d = 8'h65;	//
16'h01D3:	d = 8'h92;	//
16'h01D4:	d = 8'h44;	//
16'h01D5:	d = 8'hE2;	//
16'h01D6:	d = 8'h8F;	//
16'h01D7:	d = 8'h22;	//
16'h01D8:	d = 8'h08;	//
16'h01D9:	d = 8'h18;	//
16'h01DA:	d = 8'hC6;	//
16'h01DB:	d = 8'hE2;	//
16'h01DC:	d = 8'hF9;	//
16'h01DD:	d = 8'h23;	//
16'h01DE:	d = 8'h49;	//
16'h01DF:	d = 8'h71;	//
16'h01E0:	d = 8'h41;	//
16'h01E1:	d = 8'h20;	//
16'h01E2:	d = 8'hC3;	//
16'h01E3:	d = 8'h48;	//
16'h01E4:	d = 8'h70;	//
16'h01E5:	d = 8'h62;	//
16'h01E6:	d = 8'h7E;	//
16'h01E7:	d = 8'h0B;	//
16'h01E8:	d = 8'h1C;	//
16'h01E9:	d = 8'h0B;	//
16'h01EA:	d = 8'hA4;	//
16'h01EB:	d = 8'h35;	//
16'h01EC:	d = 8'h00;	//
16'h01ED:	d = 8'hC1;	//
16'h01EE:	d = 8'hFF;	//
16'h01EF:	d = 8'hF3;	//
16'h01F0:	d = 8'h72;	//
16'h01F1:	d = 8'h64;	//
16'h01F2:	d = 8'hF0;	//
16'h01F3:	d = 8'h14;	//
16'h01F4:	d = 8'h81;	//
16'h01F5:	d = 8'h8F;	//
16'h01F6:	d = 8'h1A;	//
16'h01F7:	d = 8'h01;	//
16'h01F8:	d = 8'h69;	//
16'h01F9:	d = 8'h89;	//
16'h01FA:	d = 8'h34;	//
16'h01FB:	d = 8'h03;	//
16'h01FC:	d = 8'h48;	//
16'h01FD:	d = 8'h03;	//
16'h01FE:	d = 8'h49;	//
16'h01FF:	d = 8'h90;	//
16'h0200:	d = 8'h2C;	//
16'h0201:	d = 8'h3B;  //
16'h0202:	d = 8'h4D;  //
16'h0203:	d = 8'hDA;  //
16'h0204:	d = 8'h25;	//
16'h0205:	d = 8'hF2;	//
16'h0206:	d = 8'hE8;	//
16'h0207:	d = 8'h21;  //
16'h0208:	d = 8'h5F;	//
16'h0209:	d = 8'hCC;	//
16'h020A:	d = 8'h88;	//
16'h020B:	d = 8'h02;	//
16'h020C:	d = 8'h37;	//
16'h020D:	d = 8'hA5;	//
16'h020E:	d = 8'h2A;	//
16'h020F:	d = 8'h92;	//
16'h0210:	d = 8'h76;	//
16'h0211:	d = 8'h45;	//
16'h0212:	d = 8'h54;	//
16'h0213:	d = 8'h66;	//
16'h0214:	d = 8'h7A;	//
16'h0215:	d = 8'h95;	//
16'h0216:	d = 8'h2B;	//
16'h0217:	d = 8'hA4;	//
16'h0218:	d = 8'h8F;	//
16'h0219:	d = 8'h66;	//
16'h021A:	d = 8'h72;	//
16'h021B:	d = 8'h5D;	//
16'h021C:	d = 8'h35;	//
16'h021D:	d = 8'h6D;	//
16'h021E:	d = 8'hE9;	//
16'h021F:	d = 8'h76;	//
16'h0220:	d = 8'hED;	//
16'h0221:	d = 8'hEB;	//
16'h0222:	d = 8'hC9;	//
16'h0223:	d = 8'hD6;	//
16'h0224:	d = 8'hAA;	//
16'h0225:	d = 8'h1B;	//
16'h0226:	d = 8'h52;	//
16'h0227:	d = 8'h26;	//
16'h0228:	d = 8'h90;	//
16'h0229:	d = 8'hC2;	//
16'h022A:	d = 8'h28;	//
16'h022B:	d = 8'hFF;	//
16'h022C:	d = 8'h10;	//
16'h022D:	d = 8'hCD;	//
16'h022E:	d = 8'h5E;	//
16'h022F:	d = 8'h5B;	//
16'h0230:	d = 8'hF4;	//
16'h0231:	d = 8'h08;	//
16'h0232:	d = 8'hF9;	//
16'h0233:	d = 8'h8C;	//
16'h0234:	d = 8'hF9;	//
16'h0235:	d = 8'hCA;	//
16'h0236:	d = 8'hCF;	//
16'h0237:	d = 8'hBC;	//
16'h0238:	d = 8'h89;	//
16'h0239:	d = 8'h38;	//
16'h023A:	d = 8'h66;	//
16'h023B:	d = 8'h93;	//
16'h023C:	d = 8'hE5;	//
16'h023D:	d = 8'hA1;	//
16'h023E:	d = 8'h91;	//
16'h023F:	d = 8'hFE;	//
16'h0240:	d = 8'hDB;	//
16'h0241:	d = 8'h35;	//
16'h0242:	d = 8'hFE;	//
16'h0243:	d = 8'h40;	//
16'h0244:	d = 8'h91;	//
16'h0245:	d = 8'h82;	//
16'h0246:	d = 8'hBB;	//
16'h0247:	d = 8'hD1;	//
16'h0248:	d = 8'hEA;	//
16'h0249:	d = 8'h41;	//
16'h024A:	d = 8'h9E;	//
16'h024B:	d = 8'hB1;	//
16'h024C:	d = 8'h1A;	//
16'h024D:	d = 8'h03;	//
16'h024E:	d = 8'h5A;	//
16'h024F:	d = 8'h38;	//
16'h0250:	d = 8'hEE;	//
16'h0251:	d = 8'h9A;	//
16'h0252:	d = 8'h2C;	//
16'h0253:	d = 8'hBA;	//
16'h0254:	d = 8'h3F;	//
16'h0255:	d = 8'h18;	//
16'h0256:	d = 8'h71;	//
16'h0257:	d = 8'hA8;	//
16'h0258:	d = 8'h73;	//
16'h0259:	d = 8'h63;	//
16'h025A:	d = 8'hC9;	//
16'h025B:	d = 8'h24;	//
16'h025C:	d = 8'hD4;	//
16'h025D:	d = 8'h5D;	//
16'h025E:	d = 8'h97;	//
16'h025F:	d = 8'hC5;	//
16'h0260:	d = 8'hB9;	//
16'h0261:	d = 8'h3F;	//
16'h0262:	d = 8'h8C;	//
16'h0263:	d = 8'hCD;	//
16'h0264:	d = 8'hFB;	//
16'h0265:	d = 8'h8A;	//
16'h0266:	d = 8'h43;	//
16'h0267:	d = 8'h2E;	//
16'h0268:	d = 8'hDB;	//
16'h0269:	d = 8'h13;	//
16'h026A:	d = 8'h8B;	//
16'h026B:	d = 8'hC0;	//
16'h026C:	d = 8'h90;	//
16'h026D:	d = 8'h3C;	//
16'h026E:	d = 8'h72;	//
16'h026F:	d = 8'h0B;	//
16'h0270:	d = 8'h8C;	//
16'h0271:	d = 8'h12;	//
16'h0272:	d = 8'hC9;	//
16'h0273:	d = 8'h74;	//
16'h0274:	d = 8'h71;	//
16'h0275:	d = 8'h79;	//
16'h0276:	d = 8'h6C;	//
16'h0277:	d = 8'hCC;	//
16'h0278:	d = 8'h13;	//
16'h0279:	d = 8'hF3;	//
16'h027A:	d = 8'h06;	//
16'h027B:	d = 8'h4E;	//
16'h027C:	d = 8'hC9;	//
16'h027D:	d = 8'h77;	//
16'h027E:	d = 8'hE6;	//
16'h027F:	d = 8'h53;	//
16'h0280:	d = 8'h16;	//
16'h0281:	d = 8'h12;	//
16'h0282:	d = 8'h05;	//
16'h0283:	d = 8'h06;	//
16'h0284:	d = 8'h25;	//
16'h0285:	d = 8'hF1;	//
16'h0286:	d = 8'hE0;	//
16'h0287:	d = 8'hF5;	//
16'h0288:	d = 8'h08;	//
16'h0289:	d = 8'hCD;	//
16'h028A:	d = 8'h7A;	//
16'h028B:	d = 8'hE7;	//
16'h028C:	d = 8'h92;	//
16'h028D:	d = 8'hAB;	//
16'h028E:	d = 8'h56;	//
16'h028F:	d = 8'h84;	//
16'h0290:	d = 8'hA1;	//
16'h0291:	d = 8'h4A;	//
16'h0292:	d = 8'h75;	//
16'h0293:	d = 8'hE1;	//
16'h0294:	d = 8'h3A;	//
16'h0295:	d = 8'h74;	//
16'h0296:	d = 8'h32;	//
16'h0297:	d = 8'hED;	//
16'h0298:	d = 8'hA6;	//
16'h0299:	d = 8'hCC;	//
16'h029A:	d = 8'h5D;	//
16'h029B:	d = 8'h59;	//
16'h029C:	d = 8'h31;	//
16'h029D:	d = 8'h11;	//
16'h029E:	d = 8'hD9;	//
16'h029F:	d = 8'hFF;	//
16'h02A0:	d = 8'hF3;	//
16'h02A1:	d = 8'h72;	//
16'h02A2:	d = 8'h64;	//
16'h02A3:	d = 8'hEE;	//
16'h02A4:	d = 8'h12;	//
16'h02A5:	d = 8'hF5;	//
16'h02A6:	d = 8'h8F;	//
16'h02A7:	d = 8'h1E;	//
16'h02A8:	d = 8'h06;	//
16'h02A9:	d = 8'h64;	//
16'h02AA:	d = 8'hC9;	//
16'h02AB:	d = 8'h7E;	//
16'h02AC:	d = 8'h03;	//
16'h02AD:	d = 8'h48;	//
16'h02AE:	d = 8'hDB;	//
16'h02AF:	d = 8'h32;	//
16'h02B0:	d = 8'hDB;	//
16'h02B1:	d = 8'hE3;	//
16'h02B2:	d = 8'h99;	//
16'h02B3:	d = 8'hFF;	//
16'h02B4:	d = 8'h2E;	//
16'h02B5:	d = 8'h43;	//
16'h02B6:	d = 8'h7C;	//
16'h02B7:	d = 8'h40;	//
16'h02B8:	d = 8'h10;	//
16'h02B9:	d = 8'h1A;	//
16'h02BA:	d = 8'h3F;	//
16'h02BB:	d = 8'hD8;	//
16'h02BC:	d = 8'h57;	//
16'h02BD:	d = 8'h96;	//
16'h02BE:	d = 8'hC9;	//
16'h02BF:	d = 8'h6B;	//
16'h02C0:	d = 8'hF9;	//
16'h02C1:	d = 8'h80;	//
16'h02C2:	d = 8'h40;	//
16'h02C3:	d = 8'h70;	//
16'h02C4:	d = 8'h71;	//
16'h02C5:	d = 8'h43;	//
16'h02C6:	d = 8'hA9;	//
16'h02C7:	d = 8'h84;	//
16'h02C8:	d = 8'h43;	//
16'h02C9:	d = 8'hD1;	//
16'h02CA:	d = 8'hEE;	//
16'h02CB:	d = 8'h33;	//
16'h02CC:	d = 8'h04;	//
16'h02CD:	d = 8'hA6;	//
16'h02CE:	d = 8'h47;	//
16'h02CF:	d = 8'h07;	//
16'h02D0:	d = 8'h31;	//
16'h02D1:	d = 8'hB1;	//
16'h02D2:	d = 8'h14;	//
16'h02D3:	d = 8'h1E;	//
16'h02D4:	d = 8'h25;	//
16'h02D5:	d = 8'hFB;	//
16'h02D6:	d = 8'h74;	//
16'h02D7:	d = 8'h51;	//
16'h02D8:	d = 8'h09;	//
16'h02D9:	d = 8'hE4;	//
16'h02DA:	d = 8'h2F;	//
16'h02DB:	d = 8'h55;	//
16'h02DC:	d = 8'hFA;	//
16'h02DD:	d = 8'h39;	//
16'h02DE:	d = 8'h75;	//
16'h02DF:	d = 8'hA9;	//
16'h02E0:	d = 8'hF1;	//
16'h02E1:	d = 8'h11;	//
16'h02E2:	d = 8'h2C;	//
16'h02E3:	d = 8'h9F;	//
16'h02E4:	d = 8'hEB;	//
16'h02E5:	d = 8'h2D;	//
16'h02E6:	d = 8'hDA;	//
16'h02E7:	d = 8'hDD;	//
16'h02E8:	d = 8'h57;	//
16'h02E9:	d = 8'h42;	//
16'h02EA:	d = 8'h5B;	//
16'h02EB:	d = 8'h6D;	//
16'h02EC:	d = 8'hC4;	//
16'h02ED:	d = 8'hC2;	//
16'h02EE:	d = 8'h41;	//
16'h02EF:	d = 8'h33;	//
16'h02F0:	d = 8'h6E;	//
16'h02F1:	d = 8'hE2;	//
16'h02F2:	d = 8'h47;	//
16'h02F3:	d = 8'h22;	//
16'h02F4:	d = 8'hA6;	//
16'h02F5:	d = 8'hAE;	//
16'h02F6:	d = 8'h2A;	//
16'h02F7:	d = 8'h09;	//
16'h02F8:	d = 8'h03;	//
16'h02F9:	d = 8'hA1;	//
16'h02FA:	d = 8'h87;	//
16'h02FB:	d = 8'h2B;	//
16'h02FC:	d = 8'h3C;	//
16'h02FD:	d = 8'h2C;	//
16'h02FE:	d = 8'h5E;	//
16'h02FF:	d = 8'h33;	//
16'h0300:	d = 8'hB7;	//
16'h0301:	d = 8'h47;  //
16'h0302:	d = 8'hC1;  //
16'h0303:	d = 8'h20;  //
16'h0304:	d = 8'h1B;	//
16'h0305:	d = 8'h83;	//
16'h0306:	d = 8'h74;	//
16'h0307:	d = 8'h69;  //
16'h0308:	d = 8'h21;	//
16'h0309:	d = 8'h1C;	//
16'h030A:	d = 8'hCB;	//
16'h030B:	d = 8'h4A;	//
16'h030C:	d = 8'h55;	//
16'h030D:	d = 8'h99;	//
16'h030E:	d = 8'hD1;	//
16'h030F:	d = 8'hD5;	//
16'h0310:	d = 8'hF4;	//
16'h0311:	d = 8'h62;	//
16'h0312:	d = 8'hAF;	//
16'h0313:	d = 8'h92;	//
16'h0314:	d = 8'h07;	//
16'h0315:	d = 8'h7F;	//
16'h0316:	d = 8'h10;	//
16'h0317:	d = 8'h48;	//
16'h0318:	d = 8'h20;	//
16'h0319:	d = 8'h28;	//
16'h031A:	d = 8'h92;	//
16'h031B:	d = 8'h7A;	//
16'h031C:	d = 8'h97;	//
16'h031D:	d = 8'h12;	//
16'h031E:	d = 8'h70;	//
16'h031F:	d = 8'hA3;	//
16'h0320:	d = 8'h29;	//
16'h0321:	d = 8'h0E;	//
16'h0322:	d = 8'h25;	//
16'h0323:	d = 8'h72;	//
16'h0324:	d = 8'hE5;	//
16'h0325:	d = 8'hE1;	//
16'h0326:	d = 8'hE8;	//
16'h0327:	d = 8'h35;	//
16'h0328:	d = 8'h2E;	//
16'h0329:	d = 8'hE9;	//
16'h032A:	d = 8'h09;	//
16'h032B:	d = 8'h6C;	//
16'h032C:	d = 8'h36;	//
16'h032D:	d = 8'h54;	//
16'h032E:	d = 8'h58;	//
16'h032F:	d = 8'h57;	//
16'h0330:	d = 8'hEE;	//
16'h0331:	d = 8'h78;	//
16'h0332:	d = 8'hAF;	//
16'h0333:	d = 8'hD4;	//
16'h0334:	d = 8'h08;	//
16'h0335:	d = 8'h5A;	//
16'h0336:	d = 8'h19;	//
16'h0337:	d = 8'h8D;	//
16'h0338:	d = 8'hC4;	//
16'h0339:	d = 8'h86;	//
16'h033A:	d = 8'hAB;	//
16'h033B:	d = 8'h9E;	//
16'h033C:	d = 8'hC9;	//
16'h033D:	d = 8'h25;	//
16'h033E:	d = 8'hEF;	//
16'h033F:	d = 8'h48;	//
16'h0340:	d = 8'h34;	//
16'h0341:	d = 8'hBB;	//
16'h0342:	d = 8'h3C;	//
16'h0343:	d = 8'h76;	//
16'h0344:	d = 8'h83;	//
16'h0345:	d = 8'h25;	//
16'h0346:	d = 8'h0A;	//
16'h0347:	d = 8'h4A;	//
16'h0348:	d = 8'h13;	//
16'h0349:	d = 8'h49;	//
16'h034A:	d = 8'hA9;	//
16'h034B:	d = 8'h6F;	//
16'h034C:	d = 8'h0A;	//
16'h034D:	d = 8'h13;	//
16'h034E:	d = 8'hFF;	//
16'h034F:	d = 8'hF3;	//
16'h0350:	d = 8'h72;	//
16'h0351:	d = 8'h64;	//
16'h0352:	d = 8'hF8;	//
16'h0353:	d = 8'h18;	//
16'h0354:	d = 8'h01;	//
16'h0355:	d = 8'h91;	//
16'h0356:	d = 8'h1E;	//
16'h0357:	d = 8'h11;	//
16'h0358:	d = 8'hAD;	//
16'h0359:	d = 8'h30;	//
16'h035A:	d = 8'h03;	//
16'h035B:	d = 8'h48;	//
16'h035C:	d = 8'h01;	//
16'h035D:	d = 8'h40;	//
16'h035E:	d = 8'hCB;	//
16'h035F:	d = 8'h4F;	//
16'h0360:	d = 8'h56;	//
16'h0361:	d = 8'h77;	//
16'h0362:	d = 8'h07;	//
16'h0363:	d = 8'h38;	//
16'h0364:	d = 8'hB3;	//
16'h0365:	d = 8'hC0;	//
16'h0366:	d = 8'hA6;	//
16'h0367:	d = 8'hDA;	//
16'h0368:	d = 8'hE2;	//
16'h0369:	d = 8'hEE;	//
16'h036A:	d = 8'h67;	//
16'h036B:	d = 8'h29;	//
16'h036C:	d = 8'hDB;	//
16'h036D:	d = 8'h61;	//
16'h036E:	d = 8'h44;	//
16'h036F:	d = 8'hD4;	//
16'h0370:	d = 8'h04;	//
16'h0371:	d = 8'h3F;	//
16'h0372:	d = 8'h0D;	//
16'h0373:	d = 8'h28;	//
16'h0374:	d = 8'hF5;	//
16'h0375:	d = 8'h56;	//
16'h0376:	d = 8'h9F;	//
16'h0377:	d = 8'hDA;	//
16'h0378:	d = 8'h3C;	//
16'h0379:	d = 8'h3F;	//
16'h037A:	d = 8'hA8;	//
16'h037B:	d = 8'h7E;	//
16'h037C:	d = 8'h58;	//
16'h037D:	d = 8'hB6;	//
16'h037E:	d = 8'hEC;	//
16'h037F:	d = 8'h6E;	//
16'h0380:	d = 8'h7E;	//
16'h0381:	d = 8'hB9;	//
16'h0382:	d = 8'h8D;	//
16'h0383:	d = 8'h46;	//
16'h0384:	d = 8'hE5;	//
16'h0385:	d = 8'h02;	//
16'h0386:	d = 8'hA6;	//
16'h0387:	d = 8'hCA;	//
16'h0388:	d = 8'h47;	//
16'h0389:	d = 8'h09;	//
16'h038A:	d = 8'hAE;	//
16'h038B:	d = 8'hCC;	//
16'h038C:	d = 8'hE5;	//
16'h038D:	d = 8'h12;	//
16'h038E:	d = 8'h1C;	//
16'h038F:	d = 8'hD5;	//
16'h0390:	d = 8'hAE;	//
16'h0391:	d = 8'h33;	//
16'h0392:	d = 8'h06;	//
16'h0393:	d = 8'h6C;	//
16'h0394:	d = 8'hE2;	//
16'h0395:	d = 8'h26;	//
16'h0396:	d = 8'hF3;	//
16'h0397:	d = 8'h35;	//
16'h0398:	d = 8'hB5;	//
16'h0399:	d = 8'hFE;	//
16'h039A:	d = 8'hA6;	//
16'h039B:	d = 8'hD5;	//
16'h039C:	d = 8'h62;	//
16'h039D:	d = 8'h6A;	//
16'h039E:	d = 8'h47;	//
16'h039F:	d = 8'hF0;	//
16'h03A0:	d = 8'hDC;	//
16'h03A1:	d = 8'h63;	//
16'h03A2:	d = 8'hE1;	//
16'h03A3:	d = 8'h4C;	//
16'h03A4:	d = 8'h94;	//
16'h03A5:	d = 8'h85;	//
16'h03A6:	d = 8'h49;	//
16'h03A7:	d = 8'hA2;	//
16'h03A8:	d = 8'h31;	//
16'h03A9:	d = 8'h6B;	//
16'h03AA:	d = 8'h35;	//
16'h03AB:	d = 8'hAE;	//
16'h03AC:	d = 8'h6B;	//
16'h03AD:	d = 8'hBC;	//
16'h03AE:	d = 8'hE6;	//
16'h03AF:	d = 8'hB4;	//
16'h03B0:	d = 8'hF7;	//
16'h03B1:	d = 8'h9B;	//
16'h03B2:	d = 8'hC3;	//
16'h03B3:	d = 8'hF1;	//
16'h03B4:	d = 8'h29;	//
16'h03B5:	d = 8'hA7;	//
16'h03B6:	d = 8'h3D;	//
16'h03B7:	d = 8'hC0;	//
16'h03B8:	d = 8'hCF;	//
16'h03B9:	d = 8'hAE;	//
16'h03BA:	d = 8'h7C;	//
16'h03BB:	d = 8'hFB;	//
16'h03BC:	d = 8'hF1;	//
16'h03BD:	d = 8'hE4;	//
16'h03BE:	d = 8'h6F;	//
16'h03BF:	d = 8'h55;	//
16'h03C0:	d = 8'hB7;	//
16'h03C1:	d = 8'h46;	//
16'h03C2:	d = 8'h6C;	//
16'h03C3:	d = 8'h8F;	//
16'h03C4:	d = 8'h0E;	//
16'h03C5:	d = 8'h9B;	//
16'h03C6:	d = 8'h92;	//
16'h03C7:	d = 8'hAC;	//
16'h03C8:	d = 8'hFE;	//
16'h03C9:	d = 8'h48;	//
16'h03CA:	d = 8'h1F;	//
16'h03CB:	d = 8'hF3;	//
16'h03CC:	d = 8'hEF;	//
16'h03CD:	d = 8'hAA;	//
16'h03CE:	d = 8'h09;	//
16'h03CF:	d = 8'h8A;	//
16'h03D0:	d = 8'h54;	//
16'h03D1:	d = 8'h60;	//
16'h03D2:	d = 8'hED;	//
16'h03D3:	d = 8'h1B;	//
16'h03D4:	d = 8'hC4;	//
16'h03D5:	d = 8'hC6;	//
16'h03D6:	d = 8'h24;	//
16'h03D7:	d = 8'hC9;	//
16'h03D8:	d = 8'hE3;	//
16'h03D9:	d = 8'hF8;	//
16'h03DA:	d = 8'h8C;	//
16'h03DB:	d = 8'hC8;	//
16'h03DC:	d = 8'h76;	//
16'h03DD:	d = 8'hB8;	//
16'h03DE:	d = 8'hAD;	//
16'h03DF:	d = 8'h44;	//
16'h03E0:	d = 8'h43;	//
16'h03E1:	d = 8'h21;	//
16'h03E2:	d = 8'h69;	//
16'h03E3:	d = 8'hC2;	//
16'h03E4:	d = 8'hD1;	//
16'h03E5:	d = 8'h66;	//
16'h03E6:	d = 8'h8F;	//
16'h03E7:	d = 8'h24;	//
16'h03E8:	d = 8'h08;	//
16'h03E9:	d = 8'h93;	//
16'h03EA:	d = 8'h45;	//
16'h03EB:	d = 8'h10;	//
16'h03EC:	d = 8'hD1;	//
16'h03ED:	d = 8'h70;	//
16'h03EE:	d = 8'hEC;	//
16'h03EF:	d = 8'h1E;	//
16'h03F0:	d = 8'hFF;	//
16'h03F1:	d = 8'hF3;	//
16'h03F2:	d = 8'h72;	//
16'h03F3:	d = 8'h64;	//
16'h03F4:	d = 8'hDA;	//
16'h03F5:	d = 8'h16;	//
16'h03F6:	d = 8'hA9;	//
16'h03F7:	d = 8'hE3;	//
16'h03F8:	d = 8'h3A;	//
16'h03F9:	d = 8'h15;	//
16'h03FA:	d = 8'hC7;	//
16'h03FB:	d = 8'hBC;	//
16'h03FC:	d = 8'h03;	//
16'h03FD:	d = 8'h48;	//
16'h03FE:	d = 8'h01;	//
16'h03FF:	d = 8'h80;	//
default:	d = 8'hFF;	//
	endcase


endmodule
