// This module receives 112 MHz as input clock
// and formes strobes for all clocked parts
// (now forms only 28 MHz strobes)

//			0       4       8       12      0       4       8       12      0       4       8       12      
//			0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 0 1 2 3 
// clk		_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-_-	112
// f0		--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__--__	56
// q0		--______--______--______--______--______--______--______--______--______--______--______--______	28
// w0		--______________--______________--______________--______________--______________--______________	14
// c0		--______________________________--______________________________--______________________________	7	(ex cbeg)
// c4		________--______________________________--______________________________--______________________	7	(ex post_cbeg)
// c8		________________--______________________________--______________________________--______________	7	(ex pre_cend)
// c12		________________________--______________________________--______________________________--______	7	(ex cend)
// c15		______________________________--______________________________--______________________________--	7


module clock (

	input wire clk,
	output reg clk175,
	output reg f0, q0, w0, c0, c4, c8, c12, c15

);


	reg [5:0] cnt = 0;

	always @(posedge clk)
		cnt <= cnt + 1;
		
		
	always @*
	begin

		f0 = cnt[0];
		q0 = cnt[1:0] == 2'd0;
		w0 = cnt[2:0] == 3'd0;
		c0 = cnt[3:0] == 4'd0;
		c4 = cnt[3:0] == 4'd4;
		c8 = cnt[3:0] == 4'd8;
		c12 = cnt[3:0] == 4'd12;
		c15 = cnt[3:0] == 4'd15;
		
		clk175 = cnt[5];
		
	end
	

endmodule
