
`include "../include/tune.v"

module rom(
	input wire [15:0] a,
	output reg [7:0] d
	
);
	
	
	always @*
	case (a)
16'h0000:	d = 8'hF3;	// di
16'h0001:	d = 8'h3C;	// inc a
16'h0002:	d = 8'hD3;	// out (0), a
16'h0003:	d = 8'h00;	// 
16'h0004:	d = 8'h18;	// jr #0001
16'h0005:	d = 8'hFB;	// 
16'h0006:	d = 8'h00;	// nop
16'h0007:	d = 8'h00;	// 
16'h0008:	d = 8'h00;	// 
16'h0009:	d = 8'h00;	// 
16'h000A:	d = 8'h00;	// 
16'h000B:	d = 8'h00;	// 
16'h000C:	d = 8'h00;	// 
16'h000D:	d = 8'h00;	// 
16'h000E:	d = 8'h00;	// 
16'h000F:	d = 8'h00;	// 
16'h0010:	d = 8'h00;	// 
16'h0011:	d = 8'h00;	// 
16'h0012:	d = 8'h00;	// 
16'h0013:	d = 8'h00;	// 
16'h0014:	d = 8'h00;	// 
16'h0015:	d = 8'h00;	// 
16'h0016:	d = 8'h00;	// 
16'h0017:	d = 8'h00;	// 
16'h0018:	d = 8'h00;	// 
16'h0019:	d = 8'h00;	// 
16'h001A:	d = 8'h00;	// 
16'h001B:	d = 8'h00;	// 
16'h001C:	d = 8'h00;	// 
16'h001D:	d = 8'h00;	// 
16'h001E:	d = 8'h00;	// 
16'h001F:	d = 8'h00;	// 
16'h0020:	d = 8'h00;	// 
16'h0021:	d = 8'h00;	// 
16'h0022:	d = 8'h00;	// 
16'h0023:	d = 8'h00;	// 
16'h0024:	d = 8'h00;	// 
16'h0025:	d = 8'h00;	// 
16'h0026:	d = 8'h00;	// 
16'h0027:	d = 8'h00;	// 
16'h0028:	d = 8'h00;	// 
16'h0029:	d = 8'h00;	// 
16'h002A:	d = 8'h00;	// 
16'h002B:	d = 8'h00;	// 
16'h002C:	d = 8'h00;	// 
16'h002D:	d = 8'h00;	// 
16'h002E:	d = 8'h00;	// 
16'h002F:	d = 8'h00;	// 
16'h0030:	d = 8'h00;	// 
16'h0031:	d = 8'h00;	// 
16'h0032:	d = 8'h00;	// 
16'h0033:	d = 8'h00;	// 
16'h0034:	d = 8'h00;	// 
16'h0035:	d = 8'h00;	// 
16'h0036:	d = 8'h00;	// 
16'h0037:	d = 8'h00;	// 
16'h0038:	d = 8'h00;	// 
16'h0039:	d = 8'h00;	// 
16'h003A:	d = 8'h00;	// 
16'h003B:	d = 8'h00;	// 
16'h003C:	d = 8'h00;	// 
16'h003D:	d = 8'h00;	// 
16'h003E:	d = 8'h00;	// 
16'h003F:	d = 8'h00;	// 
16'h0040:	d = 8'h00;	// 
16'h0041:	d = 8'h00;	// 
16'h0042:	d = 8'h00;	// 
16'h0043:	d = 8'h00;	// 
16'h0044:	d = 8'h00;	// 
16'h0045:	d = 8'h00;	// 
16'h0046:	d = 8'h00;	// 
16'h0047:	d = 8'h00;	// 
16'h0048:	d = 8'h00;	// 
16'h0049:	d = 8'h00;	// 
16'h004A:	d = 8'h00;	// 
16'h004B:	d = 8'h00;	// 
16'h004C:	d = 8'h00;	// 
16'h004D:	d = 8'h00;	// 
16'h004E:	d = 8'h00;	// 
16'h004F:	d = 8'h00;	// 
16'h0050:	d = 8'h00;	// 
16'h0051:	d = 8'h00;	// 
16'h0052:	d = 8'h00;	// 
16'h0053:	d = 8'h00;	// 
16'h0054:	d = 8'h00;	// 
16'h0055:	d = 8'h00;	// 
16'h0056:	d = 8'h00;	// 
16'h0057:	d = 8'h00;	// 
16'h0058:	d = 8'h00;	// 
16'h0059:	d = 8'h00;	// 
16'h005A:	d = 8'h00;	// 
16'h005B:	d = 8'h00;	// 
16'h005C:	d = 8'h00;	// 
16'h005D:	d = 8'h00;	// 
16'h005E:	d = 8'h00;	// 
16'h005F:	d = 8'h00;	// 
16'h0060:	d = 8'h00;	// 
16'h0061:	d = 8'h00;	// 
16'h0062:	d = 8'h00;	// 
16'h0063:	d = 8'h00;	// 
16'h0064:	d = 8'h00;	// 
16'h0065:	d = 8'h00;	// 
16'h0066:	d = 8'h00;	// 
16'h0067:	d = 8'h00;	// 
16'h0068:	d = 8'h00;	// 
16'h0069:	d = 8'h00;	// 
16'h006A:	d = 8'h00;	// 
16'h006B:	d = 8'h00;	// 
16'h006C:	d = 8'h00;	// 
16'h006D:	d = 8'h00;	// 
16'h006E:	d = 8'h00;	// 
16'h006F:	d = 8'h00;	// 
16'h0070:	d = 8'h00;	// 
16'h0071:	d = 8'h00;	// 
16'h0072:	d = 8'h00;	// 
16'h0073:	d = 8'h00;	// 
16'h0074:	d = 8'h00;	// 
16'h0075:	d = 8'h00;	// 
16'h0076:	d = 8'h00;	// 
16'h0077:	d = 8'h00;	// 
16'h0078:	d = 8'h00;	// 
16'h0079:	d = 8'h00;	// 
16'h007A:	d = 8'h00;	// 
16'h007B:	d = 8'h00;	// 
16'h007C:	d = 8'h00;	// 
16'h007D:	d = 8'h00;	// 
16'h007E:	d = 8'h00;	// 
16'h007F:	d = 8'h00;	// 
16'h0080:	d = 8'h00;	// 
16'h0081:	d = 8'h00;	// 
16'h0082:	d = 8'h00;	// 
16'h0083:	d = 8'h00;	// 
16'h0084:	d = 8'h00;	// 
16'h0085:	d = 8'h00;	// 
16'h0086:	d = 8'h00;	// 
16'h0087:	d = 8'h00;	// 
16'h0088:	d = 8'h00;	// 
16'h0089:	d = 8'h00;	// 
16'h008A:	d = 8'h00;	// 
16'h008B:	d = 8'h00;	// 
16'h008C:	d = 8'h00;	// 
16'h008D:	d = 8'h00;	// 
16'h008E:	d = 8'h00;	// 
16'h008F:	d = 8'h00;	// 
16'h0090:	d = 8'h00;	// 
16'h0091:	d = 8'h00;	// 
16'h0092:	d = 8'h00;	// 
16'h0093:	d = 8'h00;	// 
16'h0094:	d = 8'h00;	// 
16'h0095:	d = 8'h00;	// 
16'h0096:	d = 8'h00;	// 
16'h0097:	d = 8'h00;	// 
16'h0098:	d = 8'h00;	// 
16'h0099:	d = 8'h00;	// 
16'h009A:	d = 8'h00;	// 
16'h009B:	d = 8'h00;	// 
16'h009C:	d = 8'h00;	// 
16'h009D:	d = 8'h00;	// 
16'h009E:	d = 8'h00;	// 
16'h009F:	d = 8'h00;	// 
16'h00A0:	d = 8'h00;	// 
16'h00A1:	d = 8'h00;	// 
16'h00A2:	d = 8'h00;	// 
16'h00A3:	d = 8'h00;	// 
16'h00A4:	d = 8'h00;	// 
16'h00A5:	d = 8'h00;	// 
16'h00A6:	d = 8'h00;	// 
16'h00A7:	d = 8'h00;	// 
16'h00A8:	d = 8'h00;	// 
16'h00A9:	d = 8'h00;	// 
16'h00AA:	d = 8'h00;	// 
16'h00AB:	d = 8'h00;	// 
16'h00AC:	d = 8'h00;	// 
16'h00AD:	d = 8'h00;	// 
16'h00AE:	d = 8'h00;	// 
16'h00AF:	d = 8'h00;	// 
16'h00B0:	d = 8'h00;	// 
16'h00B1:	d = 8'h00;	// 
16'h00B2:	d = 8'h00;	// 
16'h00B3:	d = 8'h00;	// 
16'h00B4:	d = 8'h00;	// 
16'h00B5:	d = 8'h00;	// 
16'h00B6:	d = 8'h00;	// 
16'h00B7:	d = 8'h00;	// 
16'h00B8:	d = 8'h00;	// 
16'h00B9:	d = 8'h00;	// 
16'h00BA:	d = 8'h00;	// 
16'h00BB:	d = 8'h00;	// 
16'h00BC:	d = 8'h00;	// 
16'h00BD:	d = 8'h00;	// 
16'h00BE:	d = 8'h00;	// 
16'h00BF:	d = 8'h00;	// 
16'h00C0:	d = 8'h00;	// 
16'h00C1:	d = 8'h00;	// 
16'h00C2:	d = 8'h00;	// 
16'h00C3:	d = 8'h00;	// 
16'h00C4:	d = 8'h00;	// 
16'h00C5:	d = 8'h00;	// 
16'h00C6:	d = 8'h00;	// 
16'h00C7:	d = 8'h00;	// 
16'h00C8:	d = 8'h00;	// 
16'h00C9:	d = 8'h00;	// 
16'h00CA:	d = 8'h00;	// 
16'h00CB:	d = 8'h00;	// 
16'h00CC:	d = 8'h00;	// 
16'h00CD:	d = 8'h00;	// 
16'h00CE:	d = 8'h00;	// 
16'h00CF:	d = 8'h00;	// 
16'h00D0:	d = 8'h00;	// 
16'h00D1:	d = 8'h00;	// 
16'h00D2:	d = 8'h00;	// 
16'h00D3:	d = 8'h00;	// 
16'h00D4:	d = 8'h00;	// 
16'h00D5:	d = 8'h00;	// 
16'h00D6:	d = 8'h00;	// 
16'h00D7:	d = 8'h00;	// 
16'h00D8:	d = 8'h00;	// 
16'h00D9:	d = 8'h00;	// 
16'h00DA:	d = 8'h00;	// 
16'h00DB:	d = 8'h00;	// 
16'h00DC:	d = 8'h00;	// 
16'h00DD:	d = 8'h00;	// 
16'h00DE:	d = 8'h00;	// 
16'h00DF:	d = 8'h00;	// 
16'h00E0:	d = 8'h00;	// 
16'h00E1:	d = 8'h00;	// 
16'h00E2:	d = 8'h00;	// 
16'h00E3:	d = 8'h00;	// 
16'h00E4:	d = 8'h00;	// 
16'h00E5:	d = 8'h00;	// 
16'h00E6:	d = 8'h00;	// 
16'h00E7:	d = 8'h00;	// 
16'h00E8:	d = 8'h00;	// 
16'h00E9:	d = 8'h00;	// 
16'h00EA:	d = 8'h00;	// 
16'h00EB:	d = 8'h00;	// 
16'h00EC:	d = 8'h00;	// 
16'h00ED:	d = 8'h00;	// 
16'h00EE:	d = 8'h00;	// 
16'h00EF:	d = 8'h00;	// 
16'h00F0:	d = 8'h00;	// 
16'h00F1:	d = 8'h00;	// 
16'h00F2:	d = 8'h00;	// 
16'h00F3:	d = 8'h00;	// 
16'h00F4:	d = 8'h00;	// 
16'h00F5:	d = 8'h00;	// 
16'h00F6:	d = 8'h00;	// 
16'h00F7:	d = 8'h00;	// 
16'h00F8:	d = 8'h00;	// 
16'h00F9:	d = 8'h00;	// 
16'h00FA:	d = 8'h00;	// 
16'h00FB:	d = 8'h00;	// 
16'h00FC:	d = 8'h00;	// 
16'h00FD:	d = 8'hC3;	// 
16'h00FE:	d = 8'h00;	// 
16'h00FF:	d = 8'h00;	// 
default:	d = 8'hFF;	// 
	endcase
	
	
endmodule
